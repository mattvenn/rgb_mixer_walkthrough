magic
tech sky130A
magscale 1 2
timestamp 1647437844
<< viali >>
rect 20913 47141 20947 47175
rect 1409 47073 1443 47107
rect 3249 47073 3283 47107
rect 3985 47073 4019 47107
rect 5181 47073 5215 47107
rect 6561 47073 6595 47107
rect 8401 47073 8435 47107
rect 17417 47073 17451 47107
rect 30021 47073 30055 47107
rect 32597 47073 32631 47107
rect 36001 47073 36035 47107
rect 8953 47005 8987 47039
rect 9781 47005 9815 47039
rect 16865 47005 16899 47039
rect 20269 47005 20303 47039
rect 21097 47005 21131 47039
rect 22201 47005 22235 47039
rect 24409 47005 24443 47039
rect 27997 47005 28031 47039
rect 29561 47005 29595 47039
rect 32137 47005 32171 47039
rect 36461 47005 36495 47039
rect 37749 47005 37783 47039
rect 3065 46937 3099 46971
rect 4169 46937 4203 46971
rect 8217 46937 8251 46971
rect 17049 46937 17083 46971
rect 29745 46937 29779 46971
rect 32321 46937 32355 46971
rect 7389 46665 7423 46699
rect 7941 46597 7975 46631
rect 34437 46597 34471 46631
rect 36553 46597 36587 46631
rect 37565 46597 37599 46631
rect 4353 46529 4387 46563
rect 7481 46529 7515 46563
rect 9781 46529 9815 46563
rect 16957 46529 16991 46563
rect 20545 46529 20579 46563
rect 21189 46529 21223 46563
rect 22109 46529 22143 46563
rect 24409 46529 24443 46563
rect 27997 46529 28031 46563
rect 30481 46529 30515 46563
rect 36737 46529 36771 46563
rect 37473 46529 37507 46563
rect 1593 46461 1627 46495
rect 2053 46461 2087 46495
rect 2237 46461 2271 46495
rect 2973 46461 3007 46495
rect 4629 46461 4663 46495
rect 9597 46461 9631 46495
rect 17601 46461 17635 46495
rect 18061 46461 18095 46495
rect 18245 46461 18279 46495
rect 18705 46461 18739 46495
rect 22293 46461 22327 46495
rect 22661 46461 22695 46495
rect 24593 46461 24627 46495
rect 24869 46461 24903 46495
rect 28181 46461 28215 46495
rect 28733 46461 28767 46495
rect 32597 46461 32631 46495
rect 32781 46461 32815 46495
rect 35817 46461 35851 46495
rect 5825 46325 5859 46359
rect 6377 46325 6411 46359
rect 15025 46325 15059 46359
rect 16129 46325 16163 46359
rect 20453 46325 20487 46359
rect 21005 46325 21039 46359
rect 26985 46325 27019 46359
rect 30941 46325 30975 46359
rect 3893 46121 3927 46155
rect 4629 46121 4663 46155
rect 5181 46121 5215 46155
rect 8217 46121 8251 46155
rect 17325 46121 17359 46155
rect 18245 46121 18279 46155
rect 22569 46121 22603 46155
rect 24501 46121 24535 46155
rect 28641 46121 28675 46155
rect 29561 46121 29595 46155
rect 33333 46121 33367 46155
rect 33885 46121 33919 46155
rect 1409 45985 1443 46019
rect 5825 45985 5859 46019
rect 6469 45985 6503 46019
rect 8953 45985 8987 46019
rect 9413 45985 9447 46019
rect 14933 45985 14967 46019
rect 15485 45985 15519 46019
rect 20177 45985 20211 46019
rect 20361 45985 20395 46019
rect 21281 45985 21315 46019
rect 26249 45985 26283 46019
rect 27077 45985 27111 46019
rect 30941 45985 30975 46019
rect 31769 45985 31803 46019
rect 36277 45985 36311 46019
rect 37381 45985 37415 46019
rect 3249 45917 3283 45951
rect 3985 45917 4019 45951
rect 4721 45917 4755 45951
rect 8125 45917 8159 45951
rect 17417 45917 17451 45951
rect 18153 45917 18187 45951
rect 19441 45917 19475 45951
rect 22661 45917 22695 45951
rect 24409 45917 24443 45951
rect 28733 45917 28767 45951
rect 33241 45917 33275 45951
rect 3065 45849 3099 45883
rect 6009 45849 6043 45883
rect 9137 45849 9171 45883
rect 15117 45849 15151 45883
rect 26433 45849 26467 45883
rect 31125 45849 31159 45883
rect 36461 45849 36495 45883
rect 19349 45781 19383 45815
rect 5733 45577 5767 45611
rect 8953 45577 8987 45611
rect 25329 45577 25363 45611
rect 26341 45577 26375 45611
rect 31125 45577 31159 45611
rect 2789 45509 2823 45543
rect 15209 45509 15243 45543
rect 19165 45509 19199 45543
rect 24624 45509 24658 45543
rect 29285 45509 29319 45543
rect 32229 45509 32263 45543
rect 37381 45509 37415 45543
rect 2881 45441 2915 45475
rect 3341 45441 3375 45475
rect 5641 45441 5675 45475
rect 6561 45441 6595 45475
rect 8861 45441 8895 45475
rect 15301 45441 15335 45475
rect 20076 45441 20110 45475
rect 22385 45441 22419 45475
rect 22661 45441 22695 45475
rect 24869 45441 24903 45475
rect 25513 45441 25547 45475
rect 26249 45441 26283 45475
rect 28098 45441 28132 45475
rect 29193 45441 29227 45475
rect 31033 45441 31067 45475
rect 32137 45441 32171 45475
rect 37289 45441 37323 45475
rect 37933 45441 37967 45475
rect 1409 45373 1443 45407
rect 1685 45373 1719 45407
rect 6745 45373 6779 45407
rect 8125 45373 8159 45407
rect 17969 45373 18003 45407
rect 19349 45373 19383 45407
rect 19809 45373 19843 45407
rect 22569 45373 22603 45407
rect 28365 45373 28399 45407
rect 35817 45373 35851 45407
rect 36553 45373 36587 45407
rect 36737 45373 36771 45407
rect 23489 45305 23523 45339
rect 21189 45237 21223 45271
rect 22201 45237 22235 45271
rect 22385 45237 22419 45271
rect 26985 45237 27019 45271
rect 38025 45237 38059 45271
rect 1777 45033 1811 45067
rect 6653 45033 6687 45067
rect 7389 45033 7423 45067
rect 2329 44965 2363 44999
rect 26709 44965 26743 44999
rect 20821 44897 20855 44931
rect 23213 44897 23247 44931
rect 24409 44897 24443 44931
rect 25329 44897 25363 44931
rect 27537 44897 27571 44931
rect 37105 44897 37139 44931
rect 37933 44897 37967 44931
rect 38117 44897 38151 44931
rect 2421 44829 2455 44863
rect 6561 44829 6595 44863
rect 19533 44829 19567 44863
rect 19717 44829 19751 44863
rect 23857 44829 23891 44863
rect 24593 44829 24627 44863
rect 27353 44829 27387 44863
rect 21088 44761 21122 44795
rect 22661 44761 22695 44795
rect 22937 44761 22971 44795
rect 24777 44761 24811 44795
rect 25596 44761 25630 44795
rect 19901 44693 19935 44727
rect 22201 44693 22235 44727
rect 22845 44693 22879 44727
rect 23029 44693 23063 44727
rect 23673 44693 23707 44727
rect 27169 44693 27203 44727
rect 20177 44489 20211 44523
rect 21189 44489 21223 44523
rect 22201 44489 22235 44523
rect 27169 44489 27203 44523
rect 37473 44489 37507 44523
rect 23336 44421 23370 44455
rect 18153 44353 18187 44387
rect 18420 44353 18454 44387
rect 19993 44353 20027 44387
rect 20913 44353 20947 44387
rect 21005 44353 21039 44387
rect 23581 44353 23615 44387
rect 26065 44353 26099 44387
rect 26985 44353 27019 44387
rect 27813 44353 27847 44387
rect 29929 44353 29963 44387
rect 36737 44353 36771 44387
rect 37381 44353 37415 44387
rect 26249 44285 26283 44319
rect 19533 44149 19567 44183
rect 25881 44149 25915 44183
rect 27997 44149 28031 44183
rect 29745 44149 29779 44183
rect 19257 43945 19291 43979
rect 22017 43945 22051 43979
rect 25789 43945 25823 43979
rect 27169 43945 27203 43979
rect 21649 43809 21683 43843
rect 38117 43809 38151 43843
rect 16497 43741 16531 43775
rect 16589 43741 16623 43775
rect 16773 43741 16807 43775
rect 17417 43741 17451 43775
rect 19441 43741 19475 43775
rect 21833 43741 21867 43775
rect 25329 43741 25363 43775
rect 25973 43741 26007 43775
rect 26893 43741 26927 43775
rect 26985 43741 27019 43775
rect 27629 43741 27663 43775
rect 29561 43741 29595 43775
rect 29828 43741 29862 43775
rect 36277 43741 36311 43775
rect 27896 43673 27930 43707
rect 36461 43673 36495 43707
rect 17233 43605 17267 43639
rect 25145 43605 25179 43639
rect 29009 43605 29043 43639
rect 30941 43605 30975 43639
rect 19441 43401 19475 43435
rect 25789 43401 25823 43435
rect 27261 43401 27295 43435
rect 27353 43401 27387 43435
rect 29929 43401 29963 43435
rect 37473 43401 37507 43435
rect 17040 43333 17074 43367
rect 19901 43333 19935 43367
rect 19165 43265 19199 43299
rect 19257 43265 19291 43299
rect 20177 43265 20211 43299
rect 22937 43265 22971 43299
rect 23949 43265 23983 43299
rect 24205 43265 24239 43299
rect 25973 43265 26007 43299
rect 27169 43265 27203 43299
rect 29561 43265 29595 43299
rect 29745 43265 29779 43299
rect 31125 43265 31159 43299
rect 36093 43265 36127 43299
rect 36553 43265 36587 43299
rect 37381 43265 37415 43299
rect 16773 43197 16807 43231
rect 20085 43197 20119 43231
rect 22661 43197 22695 43231
rect 26157 43197 26191 43231
rect 25329 43129 25363 43163
rect 26985 43129 27019 43163
rect 1593 43061 1627 43095
rect 2237 43061 2271 43095
rect 18153 43061 18187 43095
rect 19901 43061 19935 43095
rect 20361 43061 20395 43095
rect 27537 43061 27571 43095
rect 31309 43061 31343 43095
rect 35909 43061 35943 43095
rect 26249 42857 26283 42891
rect 27077 42857 27111 42891
rect 19993 42789 20027 42823
rect 1409 42721 1443 42755
rect 2789 42721 2823 42755
rect 17233 42721 17267 42755
rect 23489 42721 23523 42755
rect 24869 42721 24903 42755
rect 26893 42721 26927 42755
rect 30113 42721 30147 42755
rect 16221 42653 16255 42687
rect 16865 42653 16899 42687
rect 17049 42653 17083 42687
rect 18705 42653 18739 42687
rect 21189 42653 21223 42687
rect 21465 42653 21499 42687
rect 22477 42653 22511 42687
rect 23673 42653 23707 42687
rect 25136 42653 25170 42687
rect 27077 42653 27111 42687
rect 29745 42653 29779 42687
rect 31962 42653 31996 42687
rect 32229 42653 32263 42687
rect 36277 42653 36311 42687
rect 1593 42585 1627 42619
rect 20361 42585 20395 42619
rect 22661 42585 22695 42619
rect 26801 42585 26835 42619
rect 27905 42585 27939 42619
rect 28089 42585 28123 42619
rect 29837 42585 29871 42619
rect 36461 42585 36495 42619
rect 38117 42585 38151 42619
rect 16405 42517 16439 42551
rect 18521 42517 18555 42551
rect 20177 42517 20211 42551
rect 20269 42517 20303 42551
rect 20545 42517 20579 42551
rect 22845 42517 22879 42551
rect 23857 42517 23891 42551
rect 27261 42517 27295 42551
rect 27721 42517 27755 42551
rect 29561 42517 29595 42551
rect 29929 42517 29963 42551
rect 30849 42517 30883 42551
rect 1501 42313 1535 42347
rect 19441 42313 19475 42347
rect 23949 42313 23983 42347
rect 29377 42313 29411 42347
rect 30757 42313 30791 42347
rect 37565 42313 37599 42347
rect 22477 42245 22511 42279
rect 27261 42245 27295 42279
rect 27491 42245 27525 42279
rect 29837 42245 29871 42279
rect 1593 42177 1627 42211
rect 2053 42177 2087 42211
rect 9689 42177 9723 42211
rect 18061 42177 18095 42211
rect 18328 42177 18362 42211
rect 21014 42177 21048 42211
rect 22293 42177 22327 42211
rect 22385 42177 22419 42211
rect 22615 42177 22649 42211
rect 23765 42177 23799 42211
rect 27169 42177 27203 42211
rect 27353 42177 27387 42211
rect 29561 42177 29595 42211
rect 30389 42177 30423 42211
rect 30573 42177 30607 42211
rect 33876 42177 33910 42211
rect 36553 42177 36587 42211
rect 37473 42177 37507 42211
rect 2237 42109 2271 42143
rect 2973 42109 3007 42143
rect 10425 42109 10459 42143
rect 21281 42109 21315 42143
rect 22753 42109 22787 42143
rect 27629 42109 27663 42143
rect 29745 42109 29779 42143
rect 33609 42109 33643 42143
rect 19901 41973 19935 42007
rect 22109 41973 22143 42007
rect 26985 41973 27019 42007
rect 29653 41973 29687 42007
rect 34989 41973 35023 42007
rect 2881 41769 2915 41803
rect 18613 41769 18647 41803
rect 20913 41769 20947 41803
rect 22753 41769 22787 41803
rect 33977 41769 34011 41803
rect 10057 41633 10091 41667
rect 18245 41633 18279 41667
rect 19901 41633 19935 41667
rect 29929 41633 29963 41667
rect 37105 41633 37139 41667
rect 1409 41565 1443 41599
rect 2973 41565 3007 41599
rect 9689 41565 9723 41599
rect 16221 41565 16255 41599
rect 16488 41565 16522 41599
rect 18429 41565 18463 41599
rect 20085 41565 20119 41599
rect 20269 41565 20303 41599
rect 20729 41565 20763 41599
rect 22937 41565 22971 41599
rect 27454 41565 27488 41599
rect 27721 41565 27755 41599
rect 29009 41565 29043 41599
rect 29561 41565 29595 41599
rect 29745 41565 29779 41599
rect 30849 41565 30883 41599
rect 31493 41565 31527 41599
rect 34161 41565 34195 41599
rect 36277 41565 36311 41599
rect 30941 41497 30975 41531
rect 31677 41497 31711 41531
rect 33333 41497 33367 41531
rect 36461 41497 36495 41531
rect 1593 41429 1627 41463
rect 17601 41429 17635 41463
rect 26341 41429 26375 41463
rect 28825 41429 28859 41463
rect 10517 41225 10551 41259
rect 27169 41225 27203 41259
rect 30021 41225 30055 41259
rect 31125 41225 31159 41259
rect 34253 41225 34287 41259
rect 37473 41225 37507 41259
rect 8769 41157 8803 41191
rect 9229 41157 9263 41191
rect 28908 41157 28942 41191
rect 8401 41089 8435 41123
rect 19441 41089 19475 41123
rect 19717 41089 19751 41123
rect 22661 41089 22695 41123
rect 22917 41089 22951 41123
rect 24961 41089 24995 41123
rect 26985 41089 27019 41123
rect 30941 41089 30975 41123
rect 32680 41089 32714 41123
rect 34437 41089 34471 41123
rect 35265 41089 35299 41123
rect 37381 41089 37415 41123
rect 25145 41021 25179 41055
rect 28641 41021 28675 41055
rect 32413 41021 32447 41055
rect 34621 41021 34655 41055
rect 35081 41021 35115 41055
rect 24041 40953 24075 40987
rect 33793 40953 33827 40987
rect 24777 40885 24811 40919
rect 35449 40885 35483 40919
rect 36093 40885 36127 40919
rect 36553 40885 36587 40919
rect 21005 40681 21039 40715
rect 23489 40681 23523 40715
rect 25145 40681 25179 40715
rect 32689 40681 32723 40715
rect 34161 40681 34195 40715
rect 34897 40681 34931 40715
rect 25789 40613 25823 40647
rect 11437 40545 11471 40579
rect 19533 40545 19567 40579
rect 21649 40545 21683 40579
rect 24777 40545 24811 40579
rect 24986 40545 25020 40579
rect 34989 40545 35023 40579
rect 36277 40545 36311 40579
rect 38117 40545 38151 40579
rect 1593 40477 1627 40511
rect 9689 40477 9723 40511
rect 16497 40477 16531 40511
rect 19257 40477 19291 40511
rect 23673 40477 23707 40511
rect 23857 40477 23891 40511
rect 24501 40477 24535 40511
rect 26065 40477 26099 40511
rect 27730 40477 27764 40511
rect 27997 40477 28031 40511
rect 32873 40477 32907 40511
rect 34897 40477 34931 40511
rect 35817 40477 35851 40511
rect 21097 40409 21131 40443
rect 21916 40409 21950 40443
rect 35173 40409 35207 40443
rect 36461 40409 36495 40443
rect 16681 40341 16715 40375
rect 23029 40341 23063 40375
rect 24869 40341 24903 40375
rect 25605 40341 25639 40375
rect 26617 40341 26651 40375
rect 34713 40341 34747 40375
rect 35633 40341 35667 40375
rect 18061 40137 18095 40171
rect 19901 40137 19935 40171
rect 27353 40137 27387 40171
rect 30205 40137 30239 40171
rect 3433 40069 3467 40103
rect 10517 40069 10551 40103
rect 16926 40069 16960 40103
rect 25145 40069 25179 40103
rect 30757 40069 30791 40103
rect 1593 40001 1627 40035
rect 9781 40001 9815 40035
rect 18777 40001 18811 40035
rect 20361 40001 20395 40035
rect 20545 40001 20579 40035
rect 22109 40001 22143 40035
rect 25605 40001 25639 40035
rect 25789 40001 25823 40035
rect 26985 40001 27019 40035
rect 27169 40001 27203 40035
rect 28825 40001 28859 40035
rect 29081 40001 29115 40035
rect 31585 40001 31619 40035
rect 33250 40001 33284 40035
rect 34244 40001 34278 40035
rect 36001 40001 36035 40035
rect 37289 40001 37323 40035
rect 37381 40001 37415 40035
rect 1777 39933 1811 39967
rect 16681 39933 16715 39967
rect 18521 39933 18555 39967
rect 21833 39933 21867 39967
rect 33517 39933 33551 39967
rect 33977 39933 34011 39967
rect 36185 39933 36219 39967
rect 24869 39865 24903 39899
rect 30941 39865 30975 39899
rect 20729 39797 20763 39831
rect 24685 39797 24719 39831
rect 25789 39797 25823 39831
rect 31401 39797 31435 39831
rect 32137 39797 32171 39831
rect 35357 39797 35391 39831
rect 35817 39797 35851 39831
rect 38117 39797 38151 39831
rect 2053 39593 2087 39627
rect 16773 39593 16807 39627
rect 18153 39593 18187 39627
rect 24869 39593 24903 39627
rect 28549 39593 28583 39627
rect 31125 39593 31159 39627
rect 32413 39593 32447 39627
rect 33057 39593 33091 39627
rect 34161 39593 34195 39627
rect 35265 39525 35299 39559
rect 17141 39457 17175 39491
rect 21189 39457 21223 39491
rect 30757 39457 30791 39491
rect 36277 39457 36311 39491
rect 38117 39457 38151 39491
rect 2145 39389 2179 39423
rect 16957 39389 16991 39423
rect 17969 39389 18003 39423
rect 21925 39389 21959 39423
rect 24777 39389 24811 39423
rect 25053 39389 25087 39423
rect 25145 39389 25179 39423
rect 28365 39389 28399 39423
rect 30941 39389 30975 39423
rect 32137 39389 32171 39423
rect 32229 39389 32263 39423
rect 32873 39389 32907 39423
rect 33977 39389 34011 39423
rect 35081 39389 35115 39423
rect 20922 39321 20956 39355
rect 34897 39321 34931 39355
rect 36461 39321 36495 39355
rect 19809 39253 19843 39287
rect 21741 39253 21775 39287
rect 25329 39253 25363 39287
rect 34713 39253 34747 39287
rect 34989 39253 35023 39287
rect 18337 39049 18371 39083
rect 21005 39049 21039 39083
rect 22201 39049 22235 39083
rect 32505 39049 32539 39083
rect 37565 39049 37599 39083
rect 25881 38981 25915 39015
rect 35624 38981 35658 39015
rect 14289 38913 14323 38947
rect 16865 38913 16899 38947
rect 18521 38913 18555 38947
rect 18613 38913 18647 38947
rect 19993 38913 20027 38947
rect 20177 38913 20211 38947
rect 20821 38913 20855 38947
rect 22017 38913 22051 38947
rect 24777 38913 24811 38947
rect 25053 38913 25087 38947
rect 25145 38913 25179 38947
rect 25329 38913 25363 38947
rect 25789 38913 25823 38947
rect 26065 38913 26099 38947
rect 30205 38913 30239 38947
rect 30472 38913 30506 38947
rect 32321 38913 32355 38947
rect 35357 38913 35391 38947
rect 37473 38913 37507 38947
rect 1869 38845 1903 38879
rect 2053 38845 2087 38879
rect 2881 38845 2915 38879
rect 14473 38845 14507 38879
rect 17049 38845 17083 38879
rect 21833 38845 21867 38879
rect 24961 38845 24995 38879
rect 32137 38845 32171 38879
rect 14105 38709 14139 38743
rect 16681 38709 16715 38743
rect 20361 38709 20395 38743
rect 24593 38709 24627 38743
rect 26249 38709 26283 38743
rect 31585 38709 31619 38743
rect 36737 38709 36771 38743
rect 1869 38505 1903 38539
rect 2789 38505 2823 38539
rect 17601 38505 17635 38539
rect 19901 38505 19935 38539
rect 20361 38505 20395 38539
rect 32321 38505 32355 38539
rect 18061 38437 18095 38471
rect 17785 38369 17819 38403
rect 20269 38369 20303 38403
rect 22293 38369 22327 38403
rect 32413 38369 32447 38403
rect 37105 38369 37139 38403
rect 38117 38369 38151 38403
rect 2881 38301 2915 38335
rect 15485 38301 15519 38335
rect 17877 38301 17911 38335
rect 20085 38301 20119 38335
rect 20821 38301 20855 38335
rect 21005 38301 21039 38335
rect 24593 38301 24627 38335
rect 24685 38301 24719 38335
rect 24869 38301 24903 38335
rect 24961 38301 24995 38335
rect 27445 38301 27479 38335
rect 32597 38301 32631 38335
rect 33609 38301 33643 38335
rect 35449 38301 35483 38335
rect 35633 38301 35667 38335
rect 15752 38233 15786 38267
rect 17601 38233 17635 38267
rect 20361 38233 20395 38267
rect 22560 38233 22594 38267
rect 27712 38233 27746 38267
rect 32321 38233 32355 38267
rect 33425 38233 33459 38267
rect 37933 38233 37967 38267
rect 16865 38165 16899 38199
rect 21189 38165 21223 38199
rect 23673 38165 23707 38199
rect 24409 38165 24443 38199
rect 28825 38165 28859 38199
rect 32781 38165 32815 38199
rect 33241 38165 33275 38199
rect 35817 38165 35851 38199
rect 15945 37961 15979 37995
rect 18061 37961 18095 37995
rect 20269 37961 20303 37995
rect 27629 37961 27663 37995
rect 29285 37961 29319 37995
rect 29837 37961 29871 37995
rect 32505 37961 32539 37995
rect 37473 37961 37507 37995
rect 20453 37893 20487 37927
rect 24869 37893 24903 37927
rect 26065 37893 26099 37927
rect 26249 37893 26283 37927
rect 32597 37893 32631 37927
rect 14105 37825 14139 37859
rect 16129 37825 16163 37859
rect 16937 37825 16971 37859
rect 18705 37825 18739 37859
rect 18797 37825 18831 37859
rect 19533 37825 19567 37859
rect 20085 37825 20119 37859
rect 20361 37825 20395 37859
rect 21097 37825 21131 37859
rect 23121 37825 23155 37859
rect 23305 37825 23339 37859
rect 23949 37825 23983 37859
rect 24133 37825 24167 37859
rect 24225 37825 24259 37859
rect 26985 37825 27019 37859
rect 27169 37825 27203 37859
rect 27261 37825 27295 37859
rect 27353 37825 27387 37859
rect 28917 37825 28951 37859
rect 29745 37825 29779 37859
rect 30021 37825 30055 37859
rect 32689 37825 32723 37859
rect 34529 37825 34563 37859
rect 35624 37825 35658 37859
rect 37381 37825 37415 37859
rect 16681 37757 16715 37791
rect 26433 37757 26467 37791
rect 29009 37757 29043 37791
rect 32321 37757 32355 37791
rect 35357 37757 35391 37791
rect 14289 37621 14323 37655
rect 18521 37621 18555 37655
rect 19349 37621 19383 37655
rect 20637 37621 20671 37655
rect 21281 37621 21315 37655
rect 23305 37621 23339 37655
rect 23765 37621 23799 37655
rect 24777 37621 24811 37655
rect 30021 37621 30055 37655
rect 32873 37621 32907 37655
rect 34345 37621 34379 37655
rect 36737 37621 36771 37655
rect 16773 37417 16807 37451
rect 23029 37417 23063 37451
rect 24593 37417 24627 37451
rect 27261 37417 27295 37451
rect 29009 37417 29043 37451
rect 34713 37417 34747 37451
rect 35633 37417 35667 37451
rect 17509 37349 17543 37383
rect 26249 37349 26283 37383
rect 18061 37281 18095 37315
rect 26985 37281 27019 37315
rect 27813 37281 27847 37315
rect 28549 37281 28583 37315
rect 32045 37281 32079 37315
rect 33241 37281 33275 37315
rect 35081 37281 35115 37315
rect 38117 37281 38151 37315
rect 14381 37213 14415 37247
rect 16957 37213 16991 37247
rect 19441 37213 19475 37247
rect 19625 37213 19659 37247
rect 21925 37213 21959 37247
rect 22385 37213 22419 37247
rect 22569 37213 22603 37247
rect 22664 37213 22698 37247
rect 22753 37213 22787 37247
rect 23857 37213 23891 37247
rect 24409 37213 24443 37247
rect 24593 37213 24627 37247
rect 25421 37213 25455 37247
rect 26065 37213 26099 37247
rect 26249 37213 26283 37247
rect 26893 37213 26927 37247
rect 27721 37213 27755 37247
rect 27905 37213 27939 37247
rect 28641 37213 28675 37247
rect 29561 37213 29595 37247
rect 31861 37213 31895 37247
rect 32781 37213 32815 37247
rect 33103 37213 33137 37247
rect 34897 37213 34931 37247
rect 35817 37213 35851 37247
rect 36277 37213 36311 37247
rect 14648 37145 14682 37179
rect 17693 37145 17727 37179
rect 17785 37145 17819 37179
rect 19257 37145 19291 37179
rect 21658 37145 21692 37179
rect 23673 37145 23707 37179
rect 29828 37145 29862 37179
rect 32873 37145 32907 37179
rect 32965 37145 32999 37179
rect 36461 37145 36495 37179
rect 15761 37077 15795 37111
rect 17877 37077 17911 37111
rect 20545 37077 20579 37111
rect 23489 37077 23523 37111
rect 25329 37077 25363 37111
rect 30941 37077 30975 37111
rect 31677 37077 31711 37111
rect 32597 37077 32631 37111
rect 19993 36873 20027 36907
rect 22661 36873 22695 36907
rect 23029 36873 23063 36907
rect 27169 36873 27203 36907
rect 27537 36873 27571 36907
rect 30021 36873 30055 36907
rect 32137 36873 32171 36907
rect 37473 36873 37507 36907
rect 14289 36805 14323 36839
rect 20729 36805 20763 36839
rect 20939 36805 20973 36839
rect 26065 36805 26099 36839
rect 31125 36805 31159 36839
rect 31309 36805 31343 36839
rect 34244 36805 34278 36839
rect 18613 36737 18647 36771
rect 18880 36737 18914 36771
rect 20637 36737 20671 36771
rect 20821 36737 20855 36771
rect 22845 36737 22879 36771
rect 23121 36737 23155 36771
rect 23581 36737 23615 36771
rect 23765 36737 23799 36771
rect 25329 36737 25363 36771
rect 27077 36737 27111 36771
rect 27353 36737 27387 36771
rect 29745 36737 29779 36771
rect 33250 36737 33284 36771
rect 36553 36737 36587 36771
rect 37381 36737 37415 36771
rect 15945 36669 15979 36703
rect 16129 36669 16163 36703
rect 21097 36669 21131 36703
rect 23673 36669 23707 36703
rect 30021 36669 30055 36703
rect 33517 36669 33551 36703
rect 33977 36669 34011 36703
rect 26249 36601 26283 36635
rect 29837 36601 29871 36635
rect 20453 36533 20487 36567
rect 25421 36533 25455 36567
rect 35357 36533 35391 36567
rect 14381 36329 14415 36363
rect 20269 36329 20303 36363
rect 21741 36261 21775 36295
rect 24685 36261 24719 36295
rect 26985 36261 27019 36295
rect 31585 36261 31619 36295
rect 1409 36125 1443 36159
rect 3249 36125 3283 36159
rect 14289 36125 14323 36159
rect 20361 36125 20395 36159
rect 21557 36125 21591 36159
rect 24409 36125 24443 36159
rect 25881 36125 25915 36159
rect 26065 36125 26099 36159
rect 27169 36125 27203 36159
rect 27353 36125 27387 36159
rect 31401 36125 31435 36159
rect 36277 36125 36311 36159
rect 3065 36057 3099 36091
rect 24685 36057 24719 36091
rect 36522 36057 36556 36091
rect 24501 35989 24535 36023
rect 37657 35989 37691 36023
rect 2789 35785 2823 35819
rect 36185 35785 36219 35819
rect 20168 35717 20202 35751
rect 23305 35717 23339 35751
rect 27445 35717 27479 35751
rect 2881 35649 2915 35683
rect 17417 35649 17451 35683
rect 23121 35649 23155 35683
rect 24777 35649 24811 35683
rect 24961 35649 24995 35683
rect 25513 35649 25547 35683
rect 25697 35649 25731 35683
rect 27629 35649 27663 35683
rect 33425 35649 33459 35683
rect 33885 35649 33919 35683
rect 34069 35649 34103 35683
rect 34713 35649 34747 35683
rect 36001 35649 36035 35683
rect 37841 35649 37875 35683
rect 2145 35581 2179 35615
rect 19901 35581 19935 35615
rect 24685 35581 24719 35615
rect 24869 35581 24903 35615
rect 25605 35581 25639 35615
rect 34253 35581 34287 35615
rect 38117 35581 38151 35615
rect 17233 35445 17267 35479
rect 21281 35445 21315 35479
rect 23489 35445 23523 35479
rect 24501 35445 24535 35479
rect 33241 35445 33275 35479
rect 34897 35445 34931 35479
rect 17417 35241 17451 35275
rect 20821 35241 20855 35275
rect 27721 35241 27755 35275
rect 36553 35241 36587 35275
rect 24593 35173 24627 35207
rect 26709 35173 26743 35207
rect 36093 35173 36127 35207
rect 22661 35105 22695 35139
rect 22937 35105 22971 35139
rect 24869 35105 24903 35139
rect 25789 35105 25823 35139
rect 25973 35105 26007 35139
rect 27169 35105 27203 35139
rect 27905 35105 27939 35139
rect 30021 35105 30055 35139
rect 30205 35105 30239 35139
rect 36921 35105 36955 35139
rect 15577 35037 15611 35071
rect 17601 35037 17635 35071
rect 17693 35037 17727 35071
rect 18337 35037 18371 35071
rect 18429 35037 18463 35071
rect 20637 35037 20671 35071
rect 22569 35037 22603 35071
rect 23581 35037 23615 35071
rect 23765 35037 23799 35071
rect 23857 35037 23891 35071
rect 24961 35037 24995 35071
rect 25697 35037 25731 35071
rect 25881 35037 25915 35071
rect 27077 35037 27111 35071
rect 27997 35037 28031 35071
rect 28089 35037 28123 35071
rect 28181 35037 28215 35071
rect 29929 35037 29963 35071
rect 32781 35037 32815 35071
rect 34713 35037 34747 35071
rect 36737 35037 36771 35071
rect 37473 35037 37507 35071
rect 37565 35037 37599 35071
rect 15844 34969 15878 35003
rect 31861 34969 31895 35003
rect 33048 34969 33082 35003
rect 34958 34969 34992 35003
rect 16957 34901 16991 34935
rect 18613 34901 18647 34935
rect 23397 34901 23431 34935
rect 26157 34901 26191 34935
rect 30205 34901 30239 34935
rect 31953 34901 31987 34935
rect 34161 34901 34195 34935
rect 37749 34901 37783 34935
rect 15945 34697 15979 34731
rect 18337 34697 18371 34731
rect 20821 34697 20855 34731
rect 23673 34697 23707 34731
rect 30021 34697 30055 34731
rect 33517 34697 33551 34731
rect 36185 34697 36219 34731
rect 37381 34697 37415 34731
rect 17224 34629 17258 34663
rect 32404 34629 32438 34663
rect 35725 34629 35759 34663
rect 36337 34629 36371 34663
rect 36553 34629 36587 34663
rect 16129 34561 16163 34595
rect 19910 34561 19944 34595
rect 21005 34561 21039 34595
rect 21189 34561 21223 34595
rect 22385 34561 22419 34595
rect 22564 34567 22598 34601
rect 22664 34564 22698 34598
rect 22753 34561 22787 34595
rect 23489 34561 23523 34595
rect 23673 34561 23707 34595
rect 24501 34561 24535 34595
rect 24685 34561 24719 34595
rect 24777 34561 24811 34595
rect 25053 34561 25087 34595
rect 26249 34561 26283 34595
rect 26433 34561 26467 34595
rect 27169 34561 27203 34595
rect 27353 34561 27387 34595
rect 27445 34561 27479 34595
rect 28365 34561 28399 34595
rect 29193 34561 29227 34595
rect 31134 34561 31168 34595
rect 34253 34561 34287 34595
rect 35449 34561 35483 34595
rect 37565 34561 37599 34595
rect 16957 34493 16991 34527
rect 20177 34493 20211 34527
rect 23029 34493 23063 34527
rect 24869 34493 24903 34527
rect 26341 34493 26375 34527
rect 27905 34493 27939 34527
rect 28273 34493 28307 34527
rect 28549 34493 28583 34527
rect 29285 34493 29319 34527
rect 29561 34493 29595 34527
rect 31401 34493 31435 34527
rect 32137 34493 32171 34527
rect 33977 34493 34011 34527
rect 35633 34493 35667 34527
rect 18797 34357 18831 34391
rect 25237 34357 25271 34391
rect 26985 34357 27019 34391
rect 35265 34357 35299 34391
rect 35725 34357 35759 34391
rect 36369 34357 36403 34391
rect 16681 34153 16715 34187
rect 19441 34153 19475 34187
rect 24869 34153 24903 34187
rect 27905 34153 27939 34187
rect 30573 34153 30607 34187
rect 34713 34153 34747 34187
rect 35725 34153 35759 34187
rect 16221 34085 16255 34119
rect 17877 34085 17911 34119
rect 30113 34085 30147 34119
rect 24409 34017 24443 34051
rect 29653 34017 29687 34051
rect 32137 34017 32171 34051
rect 33793 34017 33827 34051
rect 34069 34017 34103 34051
rect 34161 34017 34195 34051
rect 36737 34017 36771 34051
rect 14841 33949 14875 33983
rect 16865 33949 16899 33983
rect 17049 33949 17083 33983
rect 18153 33949 18187 33983
rect 18245 33949 18279 33983
rect 19257 33949 19291 33983
rect 21373 33949 21407 33983
rect 24501 33949 24535 33983
rect 24685 33949 24719 33983
rect 26709 33949 26743 33983
rect 26893 33949 26927 33983
rect 26985 33949 27019 33983
rect 27123 33949 27157 33983
rect 28089 33949 28123 33983
rect 28273 33949 28307 33983
rect 28365 33949 28399 33983
rect 29745 33949 29779 33983
rect 30573 33949 30607 33983
rect 30849 33949 30883 33983
rect 32413 33949 32447 33983
rect 33701 33949 33735 33983
rect 34897 33949 34931 33983
rect 34989 33949 35023 33983
rect 35909 33949 35943 33983
rect 36093 33949 36127 33983
rect 15108 33881 15142 33915
rect 21106 33881 21140 33915
rect 36001 33881 36035 33915
rect 36277 33881 36311 33915
rect 37004 33881 37038 33915
rect 18061 33813 18095 33847
rect 18429 33813 18463 33847
rect 19993 33813 20027 33847
rect 27353 33813 27387 33847
rect 30757 33813 30791 33847
rect 33517 33813 33551 33847
rect 33977 33813 34011 33847
rect 38117 33813 38151 33847
rect 15209 33609 15243 33643
rect 17785 33609 17819 33643
rect 27169 33609 27203 33643
rect 30573 33609 30607 33643
rect 34253 33609 34287 33643
rect 18245 33541 18279 33575
rect 27537 33541 27571 33575
rect 29653 33541 29687 33575
rect 15393 33473 15427 33507
rect 17969 33473 18003 33507
rect 21005 33473 21039 33507
rect 21833 33473 21867 33507
rect 25053 33473 25087 33507
rect 25320 33473 25354 33507
rect 27353 33473 27387 33507
rect 30389 33473 30423 33507
rect 34437 33473 34471 33507
rect 34713 33473 34747 33507
rect 36645 33473 36679 33507
rect 37473 33473 37507 33507
rect 37565 33473 37599 33507
rect 37749 33473 37783 33507
rect 18153 33405 18187 33439
rect 21189 33337 21223 33371
rect 34621 33337 34655 33371
rect 37289 33337 37323 33371
rect 18061 33269 18095 33303
rect 22017 33269 22051 33303
rect 26433 33269 26467 33303
rect 29561 33269 29595 33303
rect 36461 33269 36495 33303
rect 37473 33269 37507 33303
rect 15393 33065 15427 33099
rect 17325 33065 17359 33099
rect 33057 33065 33091 33099
rect 37565 33065 37599 33099
rect 30205 32929 30239 32963
rect 34713 32929 34747 32963
rect 34989 32929 35023 32963
rect 36185 32929 36219 32963
rect 15577 32861 15611 32895
rect 15669 32861 15703 32895
rect 17509 32861 17543 32895
rect 17969 32861 18003 32895
rect 23765 32861 23799 32895
rect 30481 32861 30515 32895
rect 32045 32861 32079 32895
rect 32229 32861 32263 32895
rect 32413 32861 32447 32895
rect 32873 32861 32907 32895
rect 36452 32861 36486 32895
rect 18153 32793 18187 32827
rect 18337 32725 18371 32759
rect 23673 32725 23707 32759
rect 15669 32521 15703 32555
rect 16957 32521 16991 32555
rect 23489 32521 23523 32555
rect 24317 32521 24351 32555
rect 30665 32521 30699 32555
rect 37289 32521 37323 32555
rect 28181 32453 28215 32487
rect 30297 32453 30331 32487
rect 30497 32453 30531 32487
rect 31309 32453 31343 32487
rect 32321 32453 32355 32487
rect 33324 32453 33358 32487
rect 14289 32385 14323 32419
rect 14556 32385 14590 32419
rect 16865 32385 16899 32419
rect 17049 32385 17083 32419
rect 18245 32385 18279 32419
rect 18501 32385 18535 32419
rect 20453 32385 20487 32419
rect 22109 32385 22143 32419
rect 22376 32385 22410 32419
rect 24133 32385 24167 32419
rect 24409 32385 24443 32419
rect 25329 32385 25363 32419
rect 25421 32385 25455 32419
rect 25605 32385 25639 32419
rect 27997 32385 28031 32419
rect 28273 32385 28307 32419
rect 28365 32385 28399 32419
rect 31493 32385 31527 32419
rect 32505 32385 32539 32419
rect 35265 32385 35299 32419
rect 35909 32385 35943 32419
rect 36093 32385 36127 32419
rect 36277 32385 36311 32419
rect 37473 32385 37507 32419
rect 37657 32385 37691 32419
rect 20637 32317 20671 32351
rect 33057 32317 33091 32351
rect 16681 32249 16715 32283
rect 19625 32249 19659 32283
rect 17233 32181 17267 32215
rect 20269 32181 20303 32215
rect 23949 32181 23983 32215
rect 25789 32181 25823 32215
rect 28549 32181 28583 32215
rect 30481 32181 30515 32215
rect 34437 32181 34471 32215
rect 35449 32181 35483 32215
rect 14749 31977 14783 32011
rect 16773 31977 16807 32011
rect 16957 31977 16991 32011
rect 18061 31977 18095 32011
rect 23213 31977 23247 32011
rect 26065 31977 26099 32011
rect 30941 31977 30975 32011
rect 33977 31977 34011 32011
rect 19349 31909 19383 31943
rect 20913 31909 20947 31943
rect 32045 31909 32079 31943
rect 16681 31841 16715 31875
rect 18705 31841 18739 31875
rect 20637 31841 20671 31875
rect 21097 31841 21131 31875
rect 24869 31841 24903 31875
rect 30757 31841 30791 31875
rect 36461 31841 36495 31875
rect 38117 31841 38151 31875
rect 14933 31773 14967 31807
rect 15393 31773 15427 31807
rect 15577 31773 15611 31807
rect 15761 31773 15795 31807
rect 16497 31773 16531 31807
rect 16773 31773 16807 31807
rect 18245 31773 18279 31807
rect 18337 31773 18371 31807
rect 18547 31773 18581 31807
rect 19533 31773 19567 31807
rect 22937 31773 22971 31807
rect 23029 31773 23063 31807
rect 23213 31773 23247 31807
rect 24593 31773 24627 31807
rect 24685 31773 24719 31807
rect 27353 31773 27387 31807
rect 29561 31773 29595 31807
rect 29745 31773 29779 31807
rect 29837 31773 29871 31807
rect 29929 31773 29963 31807
rect 30113 31773 30147 31807
rect 31217 31773 31251 31807
rect 32137 31773 32171 31807
rect 33057 31773 33091 31807
rect 33149 31773 33183 31807
rect 33333 31773 33367 31807
rect 33793 31773 33827 31807
rect 35817 31773 35851 31807
rect 36277 31773 36311 31807
rect 18429 31705 18463 31739
rect 24869 31637 24903 31671
rect 30297 31637 30331 31671
rect 25421 31433 25455 31467
rect 25881 31433 25915 31467
rect 30113 31433 30147 31467
rect 37565 31433 37599 31467
rect 18696 31365 18730 31399
rect 20913 31365 20947 31399
rect 21030 31365 21064 31399
rect 23020 31365 23054 31399
rect 26157 31365 26191 31399
rect 28558 31365 28592 31399
rect 29837 31365 29871 31399
rect 35602 31365 35636 31399
rect 15574 31297 15608 31331
rect 15761 31297 15795 31331
rect 16865 31297 16899 31331
rect 17049 31297 17083 31331
rect 17509 31297 17543 31331
rect 20545 31297 20579 31331
rect 24869 31297 24903 31331
rect 25145 31297 25179 31331
rect 25237 31297 25271 31331
rect 26065 31297 26099 31331
rect 26249 31297 26283 31331
rect 26433 31297 26467 31331
rect 29469 31297 29503 31331
rect 29562 31297 29596 31331
rect 29745 31297 29779 31331
rect 29975 31297 30009 31331
rect 30665 31297 30699 31331
rect 30757 31297 30791 31331
rect 32137 31297 32171 31331
rect 32404 31297 32438 31331
rect 37473 31297 37507 31331
rect 16681 31229 16715 31263
rect 18429 31229 18463 31263
rect 20821 31229 20855 31263
rect 22753 31229 22787 31263
rect 28825 31229 28859 31263
rect 35357 31229 35391 31263
rect 19809 31161 19843 31195
rect 24133 31161 24167 31195
rect 36737 31161 36771 31195
rect 15393 31093 15427 31127
rect 17693 31093 17727 31127
rect 21189 31093 21223 31127
rect 24961 31093 24995 31127
rect 27445 31093 27479 31127
rect 33517 31093 33551 31127
rect 25881 30889 25915 30923
rect 27537 30889 27571 30923
rect 28549 30889 28583 30923
rect 30389 30889 30423 30923
rect 16313 30821 16347 30855
rect 16773 30821 16807 30855
rect 20821 30821 20855 30855
rect 24593 30821 24627 30855
rect 29561 30821 29595 30855
rect 19901 30753 19935 30787
rect 21189 30753 21223 30787
rect 32413 30753 32447 30787
rect 37197 30753 37231 30787
rect 14289 30685 14323 30719
rect 14933 30685 14967 30719
rect 18153 30685 18187 30719
rect 20085 30685 20119 30719
rect 21649 30685 21683 30719
rect 21833 30685 21867 30719
rect 23029 30685 23063 30719
rect 24777 30685 24811 30719
rect 25329 30685 25363 30719
rect 25513 30685 25547 30719
rect 25697 30685 25731 30719
rect 27261 30685 27295 30719
rect 27353 30685 27387 30719
rect 27629 30685 27663 30719
rect 28089 30685 28123 30719
rect 28365 30685 28399 30719
rect 30481 30685 30515 30719
rect 31861 30685 31895 30719
rect 38117 30685 38151 30719
rect 15178 30617 15212 30651
rect 17886 30617 17920 30651
rect 20269 30617 20303 30651
rect 25605 30617 25639 30651
rect 29745 30617 29779 30651
rect 37933 30617 37967 30651
rect 14473 30549 14507 30583
rect 20729 30549 20763 30583
rect 21741 30549 21775 30583
rect 23213 30549 23247 30583
rect 27077 30549 27111 30583
rect 28181 30549 28215 30583
rect 27537 30345 27571 30379
rect 31585 30345 31619 30379
rect 37473 30345 37507 30379
rect 24961 30277 24995 30311
rect 28917 30277 28951 30311
rect 30472 30277 30506 30311
rect 33149 30277 33183 30311
rect 34336 30277 34370 30311
rect 14933 30209 14967 30243
rect 18613 30209 18647 30243
rect 20545 30209 20579 30243
rect 20729 30209 20763 30243
rect 20913 30209 20947 30243
rect 21097 30209 21131 30243
rect 22017 30209 22051 30243
rect 22109 30209 22143 30243
rect 22293 30209 22327 30243
rect 22385 30209 22419 30243
rect 24869 30209 24903 30243
rect 25053 30209 25087 30243
rect 27629 30209 27663 30243
rect 28365 30209 28399 30243
rect 28825 30209 28859 30243
rect 29469 30209 29503 30243
rect 29653 30209 29687 30243
rect 34069 30209 34103 30243
rect 37381 30209 37415 30243
rect 15393 30141 15427 30175
rect 20821 30141 20855 30175
rect 30205 30141 30239 30175
rect 28181 30073 28215 30107
rect 33425 30073 33459 30107
rect 18429 30005 18463 30039
rect 21281 30005 21315 30039
rect 21833 30005 21867 30039
rect 29469 30005 29503 30039
rect 33609 30005 33643 30039
rect 35449 30005 35483 30039
rect 36553 30005 36587 30039
rect 21097 29801 21131 29835
rect 25421 29801 25455 29835
rect 26065 29801 26099 29835
rect 26985 29801 27019 29835
rect 28825 29801 28859 29835
rect 30941 29801 30975 29835
rect 31401 29733 31435 29767
rect 32965 29733 32999 29767
rect 34161 29733 34195 29767
rect 15669 29665 15703 29699
rect 21649 29665 21683 29699
rect 28733 29665 28767 29699
rect 33517 29665 33551 29699
rect 33793 29665 33827 29699
rect 36277 29665 36311 29699
rect 38117 29665 38151 29699
rect 1777 29597 1811 29631
rect 14197 29597 14231 29631
rect 15301 29597 15335 29631
rect 20821 29597 20855 29631
rect 20913 29597 20947 29631
rect 21189 29597 21223 29631
rect 21833 29597 21867 29631
rect 22017 29597 22051 29631
rect 22109 29597 22143 29631
rect 23121 29597 23155 29631
rect 25513 29597 25547 29631
rect 25973 29597 26007 29631
rect 26893 29597 26927 29631
rect 28917 29597 28951 29631
rect 29009 29597 29043 29631
rect 29561 29597 29595 29631
rect 31677 29597 31711 29631
rect 33885 29597 33919 29631
rect 34897 29597 34931 29631
rect 34989 29597 35023 29631
rect 29806 29529 29840 29563
rect 31401 29529 31435 29563
rect 32597 29529 32631 29563
rect 34002 29529 34036 29563
rect 36461 29529 36495 29563
rect 14381 29461 14415 29495
rect 20637 29461 20671 29495
rect 23305 29461 23339 29495
rect 31585 29461 31619 29495
rect 33057 29461 33091 29495
rect 34713 29461 34747 29495
rect 24961 29257 24995 29291
rect 26985 29257 27019 29291
rect 29653 29257 29687 29291
rect 30481 29257 30515 29291
rect 37381 29257 37415 29291
rect 25145 29189 25179 29223
rect 31493 29189 31527 29223
rect 32321 29189 32355 29223
rect 33977 29189 34011 29223
rect 1685 29121 1719 29155
rect 14105 29121 14139 29155
rect 14381 29121 14415 29155
rect 14933 29121 14967 29155
rect 17969 29121 18003 29155
rect 18236 29121 18270 29155
rect 22477 29121 22511 29155
rect 22744 29121 22778 29155
rect 24869 29121 24903 29155
rect 28098 29121 28132 29155
rect 28365 29121 28399 29155
rect 29469 29121 29503 29155
rect 30665 29121 30699 29155
rect 30849 29121 30883 29155
rect 30941 29121 30975 29155
rect 31401 29119 31435 29153
rect 34437 29121 34471 29155
rect 34621 29121 34655 29155
rect 35725 29121 35759 29155
rect 37289 29121 37323 29155
rect 38117 29121 38151 29155
rect 1869 29053 1903 29087
rect 2789 29053 2823 29087
rect 15669 29053 15703 29087
rect 29285 29053 29319 29087
rect 32137 29053 32171 29087
rect 19349 28985 19383 29019
rect 23857 28985 23891 29019
rect 25145 28917 25179 28951
rect 34621 28917 34655 28951
rect 35817 28917 35851 28951
rect 36737 28917 36771 28951
rect 2237 28713 2271 28747
rect 18061 28713 18095 28747
rect 22661 28713 22695 28747
rect 25789 28713 25823 28747
rect 27629 28713 27663 28747
rect 28549 28713 28583 28747
rect 28733 28713 28767 28747
rect 17325 28577 17359 28611
rect 24409 28577 24443 28611
rect 33701 28577 33735 28611
rect 35633 28577 35667 28611
rect 35817 28577 35851 28611
rect 37105 28577 37139 28611
rect 2329 28509 2363 28543
rect 15301 28509 15335 28543
rect 18291 28509 18325 28543
rect 18426 28509 18460 28543
rect 18526 28509 18560 28543
rect 18705 28509 18739 28543
rect 22891 28509 22925 28543
rect 23029 28509 23063 28543
rect 23121 28509 23155 28543
rect 23305 28509 23339 28543
rect 26893 28509 26927 28543
rect 26985 28509 27019 28543
rect 27629 28509 27663 28543
rect 27813 28509 27847 28543
rect 33425 28509 33459 28543
rect 33609 28509 33643 28543
rect 33793 28509 33827 28543
rect 33977 28509 34011 28543
rect 34713 28509 34747 28543
rect 34989 28509 35023 28543
rect 38117 28509 38151 28543
rect 14657 28441 14691 28475
rect 17080 28441 17114 28475
rect 24676 28441 24710 28475
rect 27169 28441 27203 28475
rect 28365 28441 28399 28475
rect 15945 28373 15979 28407
rect 28565 28373 28599 28407
rect 33241 28373 33275 28407
rect 34805 28373 34839 28407
rect 35173 28373 35207 28407
rect 17325 28169 17359 28203
rect 22845 28169 22879 28203
rect 24777 28169 24811 28203
rect 25237 28169 25271 28203
rect 27261 28169 27295 28203
rect 28273 28169 28307 28203
rect 32873 28169 32907 28203
rect 19257 28101 19291 28135
rect 25605 28101 25639 28135
rect 28457 28101 28491 28135
rect 25375 28067 25409 28101
rect 12909 28033 12943 28067
rect 13645 28033 13679 28067
rect 15209 28033 15243 28067
rect 17601 28033 17635 28067
rect 17690 28033 17724 28067
rect 17790 28033 17824 28067
rect 17969 28033 18003 28067
rect 19901 28033 19935 28067
rect 20168 28033 20202 28067
rect 21833 28033 21867 28067
rect 22017 28033 22051 28067
rect 22661 28033 22695 28067
rect 22845 28033 22879 28067
rect 24777 28033 24811 28067
rect 26985 28033 27019 28067
rect 27077 28033 27111 28067
rect 28181 28033 28215 28067
rect 28917 28033 28951 28067
rect 31309 28033 31343 28067
rect 32965 28033 32999 28067
rect 33517 28033 33551 28067
rect 33793 28033 33827 28067
rect 33885 28033 33919 28067
rect 36737 28033 36771 28067
rect 37289 28033 37323 28067
rect 37933 28033 37967 28067
rect 14473 27965 14507 27999
rect 15945 27965 15979 27999
rect 24501 27965 24535 27999
rect 24685 27965 24719 27999
rect 27261 27965 27295 27999
rect 29193 27965 29227 27999
rect 33609 27965 33643 27999
rect 35725 27965 35759 27999
rect 36553 27965 36587 27999
rect 38025 27965 38059 27999
rect 13093 27897 13127 27931
rect 19441 27897 19475 27931
rect 28457 27897 28491 27931
rect 29009 27897 29043 27931
rect 31493 27897 31527 27931
rect 21281 27829 21315 27863
rect 22017 27829 22051 27863
rect 25421 27829 25455 27863
rect 29101 27829 29135 27863
rect 34069 27829 34103 27863
rect 37381 27829 37415 27863
rect 17509 27625 17543 27659
rect 20177 27625 20211 27659
rect 22293 27557 22327 27591
rect 27353 27557 27387 27591
rect 32689 27557 32723 27591
rect 15117 27489 15151 27523
rect 19349 27489 19383 27523
rect 22017 27489 22051 27523
rect 37197 27489 37231 27523
rect 37933 27489 37967 27523
rect 38117 27489 38151 27523
rect 8033 27421 8067 27455
rect 15485 27421 15519 27455
rect 16221 27421 16255 27455
rect 17417 27421 17451 27455
rect 17601 27421 17635 27455
rect 19257 27421 19291 27455
rect 19441 27421 19475 27455
rect 20453 27421 20487 27455
rect 20545 27421 20579 27455
rect 20637 27421 20671 27455
rect 20821 27421 20855 27455
rect 21925 27421 21959 27455
rect 27353 27421 27387 27455
rect 27629 27421 27663 27455
rect 30665 27421 30699 27455
rect 31309 27421 31343 27455
rect 33517 27421 33551 27455
rect 33609 27421 33643 27455
rect 33793 27421 33827 27455
rect 33885 27421 33919 27455
rect 16773 27353 16807 27387
rect 27537 27353 27571 27387
rect 31554 27353 31588 27387
rect 7849 27285 7883 27319
rect 30757 27285 30791 27319
rect 33333 27285 33367 27319
rect 17233 27081 17267 27115
rect 17785 27081 17819 27115
rect 18521 27081 18555 27115
rect 36277 27081 36311 27115
rect 8401 27013 8435 27047
rect 19165 27013 19199 27047
rect 20269 27013 20303 27047
rect 21097 27013 21131 27047
rect 29570 27013 29604 27047
rect 37841 27013 37875 27047
rect 8033 26945 8067 26979
rect 14933 26945 14967 26979
rect 16865 26945 16899 26979
rect 17877 26945 17911 26979
rect 18705 26945 18739 26979
rect 21833 26945 21867 26979
rect 21925 26945 21959 26979
rect 22109 26945 22143 26979
rect 22937 26945 22971 26979
rect 23029 26945 23063 26979
rect 23213 26945 23247 26979
rect 25145 26945 25179 26979
rect 25421 26945 25455 26979
rect 25881 26945 25915 26979
rect 25973 26945 26007 26979
rect 26157 26945 26191 26979
rect 27353 26945 27387 26979
rect 27537 26945 27571 26979
rect 30389 26945 30423 26979
rect 30573 26945 30607 26979
rect 35153 26945 35187 26979
rect 15485 26877 15519 26911
rect 16957 26877 16991 26911
rect 18797 26877 18831 26911
rect 27629 26877 27663 26911
rect 29837 26877 29871 26911
rect 34897 26877 34931 26911
rect 20453 26809 20487 26843
rect 26157 26809 26191 26843
rect 28457 26809 28491 26843
rect 21189 26741 21223 26775
rect 22293 26741 22327 26775
rect 23213 26741 23247 26775
rect 24961 26741 24995 26775
rect 25329 26741 25363 26775
rect 27169 26741 27203 26775
rect 37749 26741 37783 26775
rect 18705 26537 18739 26571
rect 21097 26537 21131 26571
rect 26065 26537 26099 26571
rect 28089 26537 28123 26571
rect 31401 26537 31435 26571
rect 34161 26537 34195 26571
rect 16405 26469 16439 26503
rect 23765 26469 23799 26503
rect 30573 26469 30607 26503
rect 16129 26401 16163 26435
rect 19533 26401 19567 26435
rect 19901 26401 19935 26435
rect 20453 26401 20487 26435
rect 20821 26401 20855 26435
rect 21557 26401 21591 26435
rect 34897 26401 34931 26435
rect 35817 26401 35851 26435
rect 36093 26401 36127 26435
rect 16037 26333 16071 26367
rect 17049 26333 17083 26367
rect 17233 26333 17267 26367
rect 17325 26333 17359 26367
rect 18337 26333 18371 26367
rect 19441 26333 19475 26367
rect 20913 26333 20947 26367
rect 22385 26333 22419 26367
rect 24685 26333 24719 26367
rect 24952 26333 24986 26367
rect 26709 26333 26743 26367
rect 30573 26333 30607 26367
rect 30849 26333 30883 26367
rect 31677 26333 31711 26367
rect 31769 26333 31803 26367
rect 31861 26333 31895 26367
rect 32045 26333 32079 26367
rect 32597 26333 32631 26367
rect 32873 26333 32907 26367
rect 33517 26333 33551 26367
rect 33701 26333 33735 26367
rect 33793 26333 33827 26367
rect 33885 26333 33919 26367
rect 34989 26333 35023 26367
rect 36185 26333 36219 26367
rect 37381 26333 37415 26367
rect 16865 26265 16899 26299
rect 18521 26265 18555 26299
rect 19257 26265 19291 26299
rect 21741 26265 21775 26299
rect 21925 26265 21959 26299
rect 22652 26265 22686 26299
rect 26976 26265 27010 26299
rect 34713 26265 34747 26299
rect 35357 26265 35391 26299
rect 37473 26265 37507 26299
rect 30757 26197 30791 26231
rect 32689 26197 32723 26231
rect 33057 26197 33091 26231
rect 17049 25993 17083 26027
rect 18613 25993 18647 26027
rect 20821 25993 20855 26027
rect 21925 25993 21959 26027
rect 22753 25993 22787 26027
rect 33241 25993 33275 26027
rect 34345 25993 34379 26027
rect 30328 25925 30362 25959
rect 31033 25925 31067 25959
rect 16129 25857 16163 25891
rect 16681 25857 16715 25891
rect 16865 25857 16899 25891
rect 18245 25857 18279 25891
rect 19257 25857 19291 25891
rect 20729 25857 20763 25891
rect 20913 25857 20947 25891
rect 21833 25857 21867 25891
rect 22017 25857 22051 25891
rect 22937 25857 22971 25891
rect 23121 25857 23155 25891
rect 25053 25857 25087 25891
rect 31217 25857 31251 25891
rect 31401 25857 31435 25891
rect 32321 25857 32355 25891
rect 33149 25857 33183 25891
rect 33333 25857 33367 25891
rect 34529 25857 34563 25891
rect 34713 25857 34747 25891
rect 35173 25857 35207 25891
rect 35357 25857 35391 25891
rect 37289 25857 37323 25891
rect 18153 25789 18187 25823
rect 19533 25789 19567 25823
rect 23213 25789 23247 25823
rect 25329 25789 25363 25823
rect 30573 25789 30607 25823
rect 31493 25789 31527 25823
rect 32229 25789 32263 25823
rect 32689 25721 32723 25755
rect 16037 25653 16071 25687
rect 19073 25653 19107 25687
rect 19441 25653 19475 25687
rect 29193 25653 29227 25687
rect 35265 25653 35299 25687
rect 36553 25653 36587 25687
rect 37381 25653 37415 25687
rect 38117 25653 38151 25687
rect 18061 25449 18095 25483
rect 25789 25449 25823 25483
rect 32229 25449 32263 25483
rect 16773 25381 16807 25415
rect 20545 25381 20579 25415
rect 18337 25313 18371 25347
rect 18429 25313 18463 25347
rect 18521 25313 18555 25347
rect 20913 25313 20947 25347
rect 24409 25313 24443 25347
rect 34989 25313 35023 25347
rect 35081 25313 35115 25347
rect 37197 25313 37231 25347
rect 37933 25313 37967 25347
rect 38117 25313 38151 25347
rect 16589 25245 16623 25279
rect 18245 25245 18279 25279
rect 19441 25245 19475 25279
rect 20729 25245 20763 25279
rect 20821 25245 20855 25279
rect 21005 25245 21039 25279
rect 30389 25245 30423 25279
rect 32045 25245 32079 25279
rect 32229 25245 32263 25279
rect 34897 25245 34931 25279
rect 35173 25245 35207 25279
rect 24654 25177 24688 25211
rect 19349 25109 19383 25143
rect 30481 25109 30515 25143
rect 34713 25109 34747 25143
rect 22033 24905 22067 24939
rect 24501 24905 24535 24939
rect 32229 24905 32263 24939
rect 34789 24905 34823 24939
rect 21833 24837 21867 24871
rect 34989 24837 35023 24871
rect 15669 24769 15703 24803
rect 15853 24769 15887 24803
rect 19717 24769 19751 24803
rect 19901 24769 19935 24803
rect 21005 24769 21039 24803
rect 21189 24769 21223 24803
rect 21281 24769 21315 24803
rect 24409 24769 24443 24803
rect 24593 24769 24627 24803
rect 27813 24769 27847 24803
rect 27905 24769 27939 24803
rect 28089 24769 28123 24803
rect 28549 24769 28583 24803
rect 32137 24769 32171 24803
rect 32321 24769 32355 24803
rect 33057 24769 33091 24803
rect 33241 24769 33275 24803
rect 33701 24769 33735 24803
rect 33885 24769 33919 24803
rect 34069 24769 34103 24803
rect 34161 24769 34195 24803
rect 35909 24769 35943 24803
rect 28641 24701 28675 24735
rect 35541 24701 35575 24735
rect 36001 24701 36035 24735
rect 34621 24633 34655 24667
rect 15761 24565 15795 24599
rect 20821 24565 20855 24599
rect 22017 24565 22051 24599
rect 22201 24565 22235 24599
rect 28089 24565 28123 24599
rect 33149 24565 33183 24599
rect 34805 24565 34839 24599
rect 37841 24565 37875 24599
rect 15761 24361 15795 24395
rect 20913 24361 20947 24395
rect 21281 24361 21315 24395
rect 35265 24361 35299 24395
rect 35633 24361 35667 24395
rect 20361 24293 20395 24327
rect 25881 24293 25915 24327
rect 26617 24293 26651 24327
rect 27353 24293 27387 24327
rect 15577 24225 15611 24259
rect 18337 24225 18371 24259
rect 22293 24225 22327 24259
rect 25697 24225 25731 24259
rect 33701 24225 33735 24259
rect 33793 24225 33827 24259
rect 36277 24225 36311 24259
rect 38117 24225 38151 24259
rect 15485 24157 15519 24191
rect 16313 24157 16347 24191
rect 16497 24157 16531 24191
rect 18245 24157 18279 24191
rect 20269 24157 20303 24191
rect 20453 24157 20487 24191
rect 21097 24157 21131 24191
rect 21373 24157 21407 24191
rect 21925 24157 21959 24191
rect 22081 24157 22115 24191
rect 22201 24157 22235 24191
rect 22477 24157 22511 24191
rect 25973 24157 26007 24191
rect 26893 24157 26927 24191
rect 28466 24157 28500 24191
rect 28733 24157 28767 24191
rect 29561 24157 29595 24191
rect 29709 24157 29743 24191
rect 29929 24157 29963 24191
rect 30026 24157 30060 24191
rect 30849 24157 30883 24191
rect 33425 24157 33459 24191
rect 33609 24157 33643 24191
rect 33977 24157 34011 24191
rect 35449 24157 35483 24191
rect 35725 24157 35759 24191
rect 26617 24089 26651 24123
rect 29837 24089 29871 24123
rect 36461 24089 36495 24123
rect 16681 24021 16715 24055
rect 18613 24021 18647 24055
rect 22661 24021 22695 24055
rect 25973 24021 26007 24055
rect 26801 24021 26835 24055
rect 30205 24021 30239 24055
rect 30757 24021 30791 24055
rect 34161 24021 34195 24055
rect 15853 23817 15887 23851
rect 15945 23817 15979 23851
rect 17693 23817 17727 23851
rect 18429 23817 18463 23851
rect 21097 23817 21131 23851
rect 22385 23817 22419 23851
rect 27721 23817 27755 23851
rect 28089 23817 28123 23851
rect 34253 23817 34287 23851
rect 36645 23817 36679 23851
rect 18337 23749 18371 23783
rect 23498 23749 23532 23783
rect 25320 23749 25354 23783
rect 32597 23749 32631 23783
rect 33425 23749 33459 23783
rect 35532 23749 35566 23783
rect 15577 23681 15611 23715
rect 16037 23681 16071 23715
rect 17325 23681 17359 23715
rect 19257 23681 19291 23715
rect 19441 23681 19475 23715
rect 20913 23681 20947 23715
rect 21097 23681 21131 23715
rect 26985 23681 27019 23715
rect 27629 23681 27663 23715
rect 27905 23681 27939 23715
rect 28549 23681 28583 23715
rect 29653 23681 29687 23715
rect 29929 23681 29963 23715
rect 30021 23681 30055 23715
rect 30205 23681 30239 23715
rect 33609 23681 33643 23715
rect 34161 23681 34195 23715
rect 34345 23681 34379 23715
rect 35265 23681 35299 23715
rect 37381 23681 37415 23715
rect 17417 23613 17451 23647
rect 18705 23613 18739 23647
rect 23765 23613 23799 23647
rect 25053 23613 25087 23647
rect 28641 23613 28675 23647
rect 29837 23613 29871 23647
rect 18613 23545 18647 23579
rect 19257 23545 19291 23579
rect 26433 23545 26467 23579
rect 27077 23545 27111 23579
rect 32781 23545 32815 23579
rect 15577 23477 15611 23511
rect 15669 23477 15703 23511
rect 18705 23477 18739 23511
rect 29469 23477 29503 23511
rect 37473 23477 37507 23511
rect 16313 23273 16347 23307
rect 19349 23273 19383 23307
rect 27077 23273 27111 23307
rect 27261 23273 27295 23307
rect 29653 23273 29687 23307
rect 15853 23205 15887 23239
rect 33793 23205 33827 23239
rect 37197 23137 37231 23171
rect 37933 23137 37967 23171
rect 38117 23137 38151 23171
rect 1777 23069 1811 23103
rect 2421 23069 2455 23103
rect 14473 23069 14507 23103
rect 14740 23069 14774 23103
rect 16313 23069 16347 23103
rect 16497 23069 16531 23103
rect 19441 23069 19475 23103
rect 21649 23069 21683 23103
rect 22109 23069 22143 23103
rect 24409 23069 24443 23103
rect 28641 23069 28675 23103
rect 28825 23069 28859 23103
rect 29009 23069 29043 23103
rect 29883 23069 29917 23103
rect 30021 23069 30055 23103
rect 30113 23069 30147 23103
rect 30297 23069 30331 23103
rect 32597 23069 32631 23103
rect 33609 23069 33643 23103
rect 35449 23069 35483 23103
rect 24676 23001 24710 23035
rect 27445 23001 27479 23035
rect 28733 23001 28767 23035
rect 32330 23001 32364 23035
rect 2329 22933 2363 22967
rect 21557 22933 21591 22967
rect 22201 22933 22235 22967
rect 25789 22933 25823 22967
rect 27235 22933 27269 22967
rect 28457 22933 28491 22967
rect 31217 22933 31251 22967
rect 35357 22933 35391 22967
rect 19257 22729 19291 22763
rect 21005 22729 21039 22763
rect 24685 22729 24719 22763
rect 32137 22729 32171 22763
rect 33885 22729 33919 22763
rect 1961 22661 1995 22695
rect 18144 22661 18178 22695
rect 22385 22661 22419 22695
rect 28825 22661 28859 22695
rect 34529 22661 34563 22695
rect 1777 22593 1811 22627
rect 16681 22593 16715 22627
rect 20637 22593 20671 22627
rect 23121 22593 23155 22627
rect 23581 22593 23615 22627
rect 23765 22593 23799 22627
rect 24593 22593 24627 22627
rect 24777 22593 24811 22627
rect 28641 22593 28675 22627
rect 29009 22593 29043 22627
rect 29469 22593 29503 22627
rect 29653 22593 29687 22627
rect 29745 22593 29779 22627
rect 30021 22593 30055 22627
rect 32413 22593 32447 22627
rect 32505 22593 32539 22627
rect 32597 22593 32631 22627
rect 32781 22593 32815 22627
rect 34989 22593 35023 22627
rect 35173 22593 35207 22627
rect 35265 22593 35299 22627
rect 35357 22593 35391 22627
rect 36277 22593 36311 22627
rect 2789 22525 2823 22559
rect 17877 22525 17911 22559
rect 20545 22525 20579 22559
rect 29837 22525 29871 22559
rect 34253 22525 34287 22559
rect 34345 22525 34379 22559
rect 36093 22525 36127 22559
rect 16773 22389 16807 22423
rect 22293 22389 22327 22423
rect 23029 22389 23063 22423
rect 23581 22389 23615 22423
rect 30205 22389 30239 22423
rect 35633 22389 35667 22423
rect 37841 22389 37875 22423
rect 26617 22185 26651 22219
rect 28273 22185 28307 22219
rect 32229 22185 32263 22219
rect 34161 22185 34195 22219
rect 20729 22117 20763 22151
rect 1869 22049 1903 22083
rect 15761 22049 15795 22083
rect 16405 22049 16439 22083
rect 16865 22049 16899 22083
rect 20453 22049 20487 22083
rect 26801 22049 26835 22083
rect 35265 22049 35299 22083
rect 35541 22049 35575 22083
rect 37197 22049 37231 22083
rect 38117 22049 38151 22083
rect 1409 21981 1443 22015
rect 15669 21981 15703 22015
rect 16589 21981 16623 22015
rect 16957 21981 16991 22015
rect 20361 21981 20395 22015
rect 22385 21981 22419 22015
rect 22477 21981 22511 22015
rect 22661 21981 22695 22015
rect 22753 21981 22787 22015
rect 23305 21981 23339 22015
rect 23397 21981 23431 22015
rect 26525 21981 26559 22015
rect 28181 21981 28215 22015
rect 32137 21981 32171 22015
rect 32321 21981 32355 22015
rect 33793 21981 33827 22015
rect 33977 21981 34011 22015
rect 35633 21981 35667 22015
rect 1593 21913 1627 21947
rect 37933 21913 37967 21947
rect 22201 21845 22235 21879
rect 26801 21845 26835 21879
rect 2053 21641 2087 21675
rect 17049 21641 17083 21675
rect 19533 21641 19567 21675
rect 20637 21641 20671 21675
rect 23121 21641 23155 21675
rect 26433 21641 26467 21675
rect 32137 21641 32171 21675
rect 34529 21641 34563 21675
rect 36461 21641 36495 21675
rect 37473 21641 37507 21675
rect 17325 21573 17359 21607
rect 17417 21573 17451 21607
rect 20913 21573 20947 21607
rect 25320 21573 25354 21607
rect 27905 21573 27939 21607
rect 29745 21573 29779 21607
rect 2145 21505 2179 21539
rect 7941 21505 7975 21539
rect 17228 21505 17262 21539
rect 17600 21505 17634 21539
rect 17693 21505 17727 21539
rect 18337 21505 18371 21539
rect 18521 21505 18555 21539
rect 18705 21505 18739 21539
rect 18889 21505 18923 21539
rect 19073 21505 19107 21539
rect 19717 21505 19751 21539
rect 19809 21505 19843 21539
rect 19901 21505 19935 21539
rect 20085 21505 20119 21539
rect 20816 21505 20850 21539
rect 21005 21505 21039 21539
rect 21188 21505 21222 21539
rect 21281 21505 21315 21539
rect 21833 21505 21867 21539
rect 22017 21505 22051 21539
rect 22385 21505 22419 21539
rect 22569 21505 22603 21539
rect 24234 21505 24268 21539
rect 24501 21505 24535 21539
rect 25053 21505 25087 21539
rect 26985 21505 27019 21539
rect 27169 21505 27203 21539
rect 27813 21505 27847 21539
rect 27997 21505 28031 21539
rect 28457 21505 28491 21539
rect 29653 21505 29687 21539
rect 30297 21505 30331 21539
rect 30481 21505 30515 21539
rect 30573 21505 30607 21539
rect 30665 21505 30699 21539
rect 32505 21505 32539 21539
rect 33149 21505 33183 21539
rect 33333 21505 33367 21539
rect 34437 21505 34471 21539
rect 34621 21505 34655 21539
rect 35081 21505 35115 21539
rect 35348 21505 35382 21539
rect 37381 21505 37415 21539
rect 8769 21437 8803 21471
rect 18797 21437 18831 21471
rect 22201 21437 22235 21471
rect 22293 21437 22327 21471
rect 32413 21437 32447 21471
rect 33241 21437 33275 21471
rect 27353 21301 27387 21335
rect 28641 21301 28675 21335
rect 30849 21301 30883 21335
rect 1685 21097 1719 21131
rect 16129 21097 16163 21131
rect 16589 21097 16623 21131
rect 19993 21097 20027 21131
rect 26525 21097 26559 21131
rect 27353 21097 27387 21131
rect 28457 21097 28491 21131
rect 31861 21097 31895 21131
rect 9873 21029 9907 21063
rect 8217 20961 8251 20995
rect 23029 20961 23063 20995
rect 23305 20961 23339 20995
rect 26709 20961 26743 20995
rect 30205 20961 30239 20995
rect 31401 20961 31435 20995
rect 31493 20961 31527 20995
rect 33609 20961 33643 20995
rect 33885 20961 33919 20995
rect 34713 20961 34747 20995
rect 38117 20961 38151 20995
rect 7941 20893 7975 20927
rect 9781 20893 9815 20927
rect 16313 20893 16347 20927
rect 16405 20893 16439 20927
rect 16681 20893 16715 20927
rect 20177 20893 20211 20927
rect 26433 20893 26467 20927
rect 28365 20893 28399 20927
rect 29929 20893 29963 20927
rect 30113 20893 30147 20927
rect 30297 20893 30331 20927
rect 30481 20893 30515 20927
rect 31125 20893 31159 20927
rect 31309 20893 31343 20927
rect 31677 20893 31711 20927
rect 32505 20893 32539 20927
rect 32689 20893 32723 20927
rect 32781 20893 32815 20927
rect 33793 20893 33827 20927
rect 33977 20893 34011 20927
rect 34069 20893 34103 20927
rect 35081 20893 35115 20927
rect 35173 20893 35207 20927
rect 36277 20893 36311 20927
rect 20361 20825 20395 20859
rect 27321 20825 27355 20859
rect 27537 20825 27571 20859
rect 30665 20825 30699 20859
rect 36461 20825 36495 20859
rect 26709 20757 26743 20791
rect 27169 20757 27203 20791
rect 32321 20757 32355 20791
rect 35357 20757 35391 20791
rect 26433 20553 26467 20587
rect 29561 20553 29595 20587
rect 33057 20553 33091 20587
rect 33701 20553 33735 20587
rect 34253 20553 34287 20587
rect 7941 20485 7975 20519
rect 15761 20485 15795 20519
rect 17785 20485 17819 20519
rect 22905 20485 22939 20519
rect 23121 20485 23155 20519
rect 23765 20485 23799 20519
rect 25320 20485 25354 20519
rect 27077 20485 27111 20519
rect 29837 20485 29871 20519
rect 15577 20417 15611 20451
rect 15853 20417 15887 20451
rect 16681 20417 16715 20451
rect 16865 20417 16899 20451
rect 17509 20417 17543 20451
rect 23581 20417 23615 20451
rect 23857 20417 23891 20451
rect 25053 20417 25087 20451
rect 26985 20417 27019 20451
rect 27169 20417 27203 20451
rect 28641 20417 28675 20451
rect 28733 20417 28767 20451
rect 29699 20417 29733 20451
rect 29929 20417 29963 20451
rect 30112 20417 30146 20451
rect 30205 20417 30239 20451
rect 30941 20417 30975 20451
rect 32689 20417 32723 20451
rect 32873 20417 32907 20451
rect 33609 20417 33643 20451
rect 34437 20417 34471 20451
rect 36553 20417 36587 20451
rect 37381 20417 37415 20451
rect 9597 20349 9631 20383
rect 17785 20349 17819 20383
rect 31033 20349 31067 20383
rect 34713 20349 34747 20383
rect 31309 20281 31343 20315
rect 34621 20281 34655 20315
rect 1593 20213 1627 20247
rect 15577 20213 15611 20247
rect 16865 20213 16899 20247
rect 17601 20213 17635 20247
rect 22753 20213 22787 20247
rect 22937 20213 22971 20247
rect 23581 20213 23615 20247
rect 37473 20213 37507 20247
rect 15577 20009 15611 20043
rect 17877 20009 17911 20043
rect 18061 20009 18095 20043
rect 19717 20009 19751 20043
rect 29745 20009 29779 20043
rect 30757 20009 30791 20043
rect 32413 20009 32447 20043
rect 21925 19941 21959 19975
rect 1409 19873 1443 19907
rect 1869 19873 1903 19907
rect 14197 19873 14231 19907
rect 20637 19873 20671 19907
rect 22569 19873 22603 19907
rect 22845 19873 22879 19907
rect 27353 19873 27387 19907
rect 37197 19873 37231 19907
rect 37933 19873 37967 19907
rect 7757 19805 7791 19839
rect 16037 19805 16071 19839
rect 20361 19805 20395 19839
rect 20453 19805 20487 19839
rect 21833 19805 21867 19839
rect 22109 19805 22143 19839
rect 25053 19805 25087 19839
rect 27537 19805 27571 19839
rect 27629 19805 27663 19839
rect 28089 19805 28123 19839
rect 28273 19805 28307 19839
rect 29653 19805 29687 19839
rect 30849 19805 30883 19839
rect 32229 19805 32263 19839
rect 32413 19805 32447 19839
rect 38117 19805 38151 19839
rect 1593 19737 1627 19771
rect 8125 19737 8159 19771
rect 14464 19737 14498 19771
rect 16304 19737 16338 19771
rect 18245 19737 18279 19771
rect 19901 19737 19935 19771
rect 24869 19737 24903 19771
rect 27353 19737 27387 19771
rect 17417 19669 17451 19703
rect 18045 19669 18079 19703
rect 19533 19669 19567 19703
rect 19701 19669 19735 19703
rect 20637 19669 20671 19703
rect 21833 19669 21867 19703
rect 28181 19669 28215 19703
rect 1961 19465 1995 19499
rect 17601 19465 17635 19499
rect 18061 19465 18095 19499
rect 19901 19465 19935 19499
rect 23213 19465 23247 19499
rect 23673 19465 23707 19499
rect 26985 19465 27019 19499
rect 29377 19465 29411 19499
rect 24786 19397 24820 19431
rect 2053 19329 2087 19363
rect 15485 19329 15519 19363
rect 15669 19329 15703 19363
rect 17417 19329 17451 19363
rect 19185 19329 19219 19363
rect 19441 19329 19475 19363
rect 21014 19329 21048 19363
rect 21281 19329 21315 19363
rect 21833 19329 21867 19363
rect 22100 19329 22134 19363
rect 25053 19329 25087 19363
rect 26249 19329 26283 19363
rect 26433 19329 26467 19363
rect 27169 19329 27203 19363
rect 27997 19329 28031 19363
rect 28264 19329 28298 19363
rect 34437 19329 34471 19363
rect 37841 19329 37875 19363
rect 15301 19261 15335 19295
rect 15761 19261 15795 19295
rect 17233 19261 17267 19295
rect 27353 19261 27387 19295
rect 34069 19261 34103 19295
rect 34345 19261 34379 19295
rect 26433 19125 26467 19159
rect 17877 18921 17911 18955
rect 19441 18921 19475 18955
rect 20913 18921 20947 18955
rect 22109 18921 22143 18955
rect 22477 18921 22511 18955
rect 27905 18921 27939 18955
rect 28089 18921 28123 18955
rect 28917 18921 28951 18955
rect 23029 18853 23063 18887
rect 29561 18853 29595 18887
rect 17969 18785 18003 18819
rect 20269 18785 20303 18819
rect 26893 18785 26927 18819
rect 31769 18785 31803 18819
rect 35173 18785 35207 18819
rect 17693 18717 17727 18751
rect 18429 18717 18463 18751
rect 18613 18717 18647 18751
rect 19257 18717 19291 18751
rect 19441 18717 19475 18751
rect 20085 18717 20119 18751
rect 20729 18717 20763 18751
rect 20913 18717 20947 18751
rect 22293 18717 22327 18751
rect 22569 18717 22603 18751
rect 23305 18717 23339 18751
rect 26617 18717 26651 18751
rect 26801 18717 26835 18751
rect 28733 18717 28767 18751
rect 29009 18717 29043 18751
rect 29837 18717 29871 18751
rect 30849 18717 30883 18751
rect 31033 18717 31067 18751
rect 31861 18717 31895 18751
rect 32873 18717 32907 18751
rect 33057 18717 33091 18751
rect 35081 18717 35115 18751
rect 36277 18717 36311 18751
rect 18521 18649 18555 18683
rect 19901 18649 19935 18683
rect 23029 18649 23063 18683
rect 27721 18649 27755 18683
rect 29561 18649 29595 18683
rect 29745 18649 29779 18683
rect 36461 18649 36495 18683
rect 38117 18649 38151 18683
rect 17509 18581 17543 18615
rect 23213 18581 23247 18615
rect 26433 18581 26467 18615
rect 27921 18581 27955 18615
rect 28549 18581 28583 18615
rect 30941 18581 30975 18615
rect 31493 18581 31527 18615
rect 32965 18581 32999 18615
rect 34713 18581 34747 18615
rect 18429 18377 18463 18411
rect 19349 18377 19383 18411
rect 29837 18377 29871 18411
rect 31493 18377 31527 18411
rect 34345 18377 34379 18411
rect 37565 18377 37599 18411
rect 17049 18241 17083 18275
rect 17316 18241 17350 18275
rect 19625 18241 19659 18275
rect 28457 18241 28491 18275
rect 28713 18241 28747 18275
rect 31309 18241 31343 18275
rect 31585 18241 31619 18275
rect 32965 18241 32999 18275
rect 33232 18241 33266 18275
rect 36553 18241 36587 18275
rect 37473 18241 37507 18275
rect 19349 18173 19383 18207
rect 19533 18173 19567 18207
rect 31217 18173 31251 18207
rect 1685 18037 1719 18071
rect 31217 18037 31251 18071
rect 36093 18037 36127 18071
rect 27169 17833 27203 17867
rect 30205 17833 30239 17867
rect 33057 17833 33091 17867
rect 32873 17765 32907 17799
rect 1409 17697 1443 17731
rect 2789 17697 2823 17731
rect 25789 17697 25823 17731
rect 31585 17697 31619 17731
rect 32965 17697 32999 17731
rect 36277 17697 36311 17731
rect 38117 17697 38151 17731
rect 26056 17629 26090 17663
rect 33149 17629 33183 17663
rect 33333 17629 33367 17663
rect 1593 17561 1627 17595
rect 31318 17561 31352 17595
rect 36461 17561 36495 17595
rect 2145 17289 2179 17323
rect 37565 17289 37599 17323
rect 2237 17153 2271 17187
rect 37473 17153 37507 17187
rect 1409 16949 1443 16983
rect 36553 16949 36587 16983
rect 1409 16609 1443 16643
rect 1869 16609 1903 16643
rect 36277 16609 36311 16643
rect 38117 16609 38151 16643
rect 1593 16473 1627 16507
rect 36461 16473 36495 16507
rect 2053 16201 2087 16235
rect 37565 16201 37599 16235
rect 2145 16065 2179 16099
rect 37473 16065 37507 16099
rect 2789 15861 2823 15895
rect 36553 15861 36587 15895
rect 1409 15521 1443 15555
rect 3249 15521 3283 15555
rect 36277 15521 36311 15555
rect 38117 15521 38151 15555
rect 3065 15385 3099 15419
rect 36461 15385 36495 15419
rect 1961 15113 1995 15147
rect 36553 15113 36587 15147
rect 1869 14977 1903 15011
rect 36461 14977 36495 15011
rect 1777 14365 1811 14399
rect 1685 13889 1719 13923
rect 1869 13821 1903 13855
rect 2789 13821 2823 13855
rect 2145 13481 2179 13515
rect 1593 13277 1627 13311
rect 2237 13277 2271 13311
rect 37841 12869 37875 12903
rect 1685 12801 1719 12835
rect 38117 12801 38151 12835
rect 1869 12733 1903 12767
rect 2789 12733 2823 12767
rect 2145 12393 2179 12427
rect 2237 12189 2271 12223
rect 37841 12189 37875 12223
rect 37381 11713 37415 11747
rect 37473 11509 37507 11543
rect 37197 11169 37231 11203
rect 37933 11169 37967 11203
rect 38117 11169 38151 11203
rect 2053 11101 2087 11135
rect 2697 11101 2731 11135
rect 1961 11033 1995 11067
rect 3249 10693 3283 10727
rect 3433 10625 3467 10659
rect 37473 10625 37507 10659
rect 1593 10557 1627 10591
rect 37381 10421 37415 10455
rect 38117 10421 38151 10455
rect 36461 10081 36495 10115
rect 1869 10013 1903 10047
rect 2513 10013 2547 10047
rect 36277 10013 36311 10047
rect 38117 9945 38151 9979
rect 2421 9877 2455 9911
rect 2053 9605 2087 9639
rect 1869 9537 1903 9571
rect 36553 9537 36587 9571
rect 37473 9537 37507 9571
rect 2789 9469 2823 9503
rect 37565 9333 37599 9367
rect 37197 8993 37231 9027
rect 37933 8993 37967 9027
rect 38117 8993 38151 9027
rect 2053 8925 2087 8959
rect 2697 8925 2731 8959
rect 2605 8789 2639 8823
rect 2237 8517 2271 8551
rect 2053 8449 2087 8483
rect 2881 8381 2915 8415
rect 37841 8313 37875 8347
rect 1409 8245 1443 8279
rect 1409 7905 1443 7939
rect 2789 7905 2823 7939
rect 37841 7837 37875 7871
rect 1593 7769 1627 7803
rect 2237 7497 2271 7531
rect 2329 7361 2363 7395
rect 37473 7361 37507 7395
rect 1501 7157 1535 7191
rect 37565 7157 37599 7191
rect 1409 6817 1443 6851
rect 2789 6817 2823 6851
rect 37197 6817 37231 6851
rect 37933 6817 37967 6851
rect 38117 6817 38151 6851
rect 1593 6681 1627 6715
rect 2053 6409 2087 6443
rect 2145 6273 2179 6307
rect 37473 6273 37507 6307
rect 35357 6205 35391 6239
rect 36553 6205 36587 6239
rect 36737 6205 36771 6239
rect 2789 6069 2823 6103
rect 37565 6069 37599 6103
rect 3249 5729 3283 5763
rect 37197 5729 37231 5763
rect 37933 5729 37967 5763
rect 38117 5729 38151 5763
rect 33425 5661 33459 5695
rect 34897 5661 34931 5695
rect 35725 5661 35759 5695
rect 1409 5593 1443 5627
rect 3065 5593 3099 5627
rect 35633 5525 35667 5559
rect 1961 5321 1995 5355
rect 36277 5321 36311 5355
rect 35265 5253 35299 5287
rect 2053 5185 2087 5219
rect 32689 5185 32723 5219
rect 33425 5185 33459 5219
rect 36369 5185 36403 5219
rect 37289 5185 37323 5219
rect 37933 5185 37967 5219
rect 2973 5117 3007 5151
rect 3157 5117 3191 5151
rect 3985 5117 4019 5151
rect 32781 5117 32815 5151
rect 33609 5117 33643 5151
rect 37381 5049 37415 5083
rect 6377 4981 6411 5015
rect 7481 4981 7515 5015
rect 2973 4777 3007 4811
rect 3893 4777 3927 4811
rect 5273 4641 5307 4675
rect 6377 4641 6411 4675
rect 6837 4641 6871 4675
rect 15669 4641 15703 4675
rect 33701 4641 33735 4675
rect 33977 4641 34011 4675
rect 34161 4641 34195 4675
rect 35541 4641 35575 4675
rect 36093 4641 36127 4675
rect 1593 4573 1627 4607
rect 3985 4573 4019 4607
rect 4629 4573 4663 4607
rect 5917 4573 5951 4607
rect 9413 4573 9447 4607
rect 9873 4573 9907 4607
rect 15209 4573 15243 4607
rect 22385 4573 22419 4607
rect 34897 4573 34931 4607
rect 35357 4573 35391 4607
rect 37657 4573 37691 4607
rect 6561 4505 6595 4539
rect 15393 4505 15427 4539
rect 9321 4437 9355 4471
rect 15577 4233 15611 4267
rect 4721 4097 4755 4131
rect 6561 4097 6595 4131
rect 7297 4097 7331 4131
rect 7389 4097 7423 4131
rect 11713 4097 11747 4131
rect 15669 4097 15703 4131
rect 20361 4097 20395 4131
rect 22201 4097 22235 4131
rect 32229 4097 32263 4131
rect 37381 4097 37415 4131
rect 1961 4029 1995 4063
rect 2145 4029 2179 4063
rect 2605 4029 2639 4063
rect 8033 4029 8067 4063
rect 8493 4029 8527 4063
rect 8677 4029 8711 4063
rect 9321 4029 9355 4063
rect 23397 4029 23431 4063
rect 23581 4029 23615 4063
rect 23857 4029 23891 4063
rect 32505 4029 32539 4063
rect 34805 4029 34839 4063
rect 34989 4029 35023 4063
rect 35449 4029 35483 4063
rect 4813 3893 4847 3927
rect 5365 3893 5399 3927
rect 6469 3893 6503 3927
rect 10793 3893 10827 3927
rect 11805 3893 11839 3927
rect 18153 3893 18187 3927
rect 20269 3893 20303 3927
rect 22293 3893 22327 3927
rect 37473 3893 37507 3927
rect 2513 3689 2547 3723
rect 9229 3689 9263 3723
rect 34161 3689 34195 3723
rect 35081 3689 35115 3723
rect 15117 3621 15151 3655
rect 22569 3621 22603 3655
rect 23121 3621 23155 3655
rect 4629 3553 4663 3587
rect 4813 3553 4847 3587
rect 5181 3553 5215 3587
rect 10425 3553 10459 3587
rect 10977 3553 11011 3587
rect 16773 3553 16807 3587
rect 20177 3553 20211 3587
rect 20637 3553 20671 3587
rect 24409 3553 24443 3587
rect 24593 3553 24627 3587
rect 24869 3553 24903 3587
rect 1961 3485 1995 3519
rect 2605 3485 2639 3519
rect 3065 3485 3099 3519
rect 3801 3485 3835 3519
rect 7113 3485 7147 3519
rect 8309 3485 8343 3519
rect 9321 3485 9355 3519
rect 9781 3485 9815 3519
rect 12725 3485 12759 3519
rect 15577 3485 15611 3519
rect 16221 3485 16255 3519
rect 18705 3485 18739 3519
rect 19533 3485 19567 3519
rect 19993 3485 20027 3519
rect 23029 3485 23063 3519
rect 23673 3485 23707 3519
rect 28181 3485 28215 3519
rect 28641 3485 28675 3519
rect 32689 3485 32723 3519
rect 33333 3485 33367 3519
rect 35173 3485 35207 3519
rect 35633 3485 35667 3519
rect 38117 3485 38151 3519
rect 9873 3417 9907 3451
rect 10609 3417 10643 3451
rect 15669 3417 15703 3451
rect 16405 3417 16439 3451
rect 36277 3417 36311 3451
rect 37933 3417 37967 3451
rect 1869 3349 1903 3383
rect 3157 3349 3191 3383
rect 7021 3349 7055 3383
rect 8217 3349 8251 3383
rect 18613 3349 18647 3383
rect 23765 3349 23799 3383
rect 28089 3349 28123 3383
rect 32781 3349 32815 3383
rect 35725 3349 35759 3383
rect 37473 3145 37507 3179
rect 3157 3077 3191 3111
rect 6837 3077 6871 3111
rect 9137 3077 9171 3111
rect 11897 3077 11931 3111
rect 18337 3077 18371 3111
rect 24041 3077 24075 3111
rect 27997 3077 28031 3111
rect 33425 3077 33459 3111
rect 1961 3009 1995 3043
rect 2973 3009 3007 3043
rect 5457 3009 5491 3043
rect 6653 3009 6687 3043
rect 8953 3009 8987 3043
rect 11713 3009 11747 3043
rect 16681 3009 16715 3043
rect 18153 3009 18187 3043
rect 27813 3009 27847 3043
rect 33241 3009 33275 3043
rect 37381 3009 37415 3043
rect 3433 2941 3467 2975
rect 7113 2941 7147 2975
rect 9413 2941 9447 2975
rect 12265 2941 12299 2975
rect 18705 2941 18739 2975
rect 23397 2941 23431 2975
rect 23857 2941 23891 2975
rect 24501 2941 24535 2975
rect 28365 2941 28399 2975
rect 35081 2941 35115 2975
rect 5365 2805 5399 2839
rect 36001 2805 36035 2839
rect 22017 2601 22051 2635
rect 37841 2601 37875 2635
rect 1409 2465 1443 2499
rect 1593 2465 1627 2499
rect 2789 2465 2823 2499
rect 5641 2465 5675 2499
rect 5825 2465 5859 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 6837 2465 6871 2499
rect 9045 2465 9079 2499
rect 9229 2465 9263 2499
rect 9689 2465 9723 2499
rect 33701 2465 33735 2499
rect 34161 2465 34195 2499
rect 34897 2465 34931 2499
rect 21833 2397 21867 2431
rect 3985 2329 4019 2363
rect 33977 2329 34011 2363
rect 35081 2329 35115 2363
rect 36737 2329 36771 2363
<< metal1 >>
rect 35894 47404 35900 47456
rect 35952 47444 35958 47456
rect 37182 47444 37188 47456
rect 35952 47416 37188 47444
rect 35952 47404 35958 47416
rect 37182 47404 37188 47416
rect 37240 47404 37246 47456
rect 1104 47354 38824 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 38824 47354
rect 1104 47280 38824 47302
rect 3326 47132 3332 47184
rect 3384 47172 3390 47184
rect 3384 47144 6592 47172
rect 3384 47132 3390 47144
rect 1394 47104 1400 47116
rect 1355 47076 1400 47104
rect 1394 47064 1400 47076
rect 1452 47064 1458 47116
rect 2866 47064 2872 47116
rect 2924 47104 2930 47116
rect 3237 47107 3295 47113
rect 3237 47104 3249 47107
rect 2924 47076 3249 47104
rect 2924 47064 2930 47076
rect 3237 47073 3249 47076
rect 3283 47073 3295 47107
rect 3237 47067 3295 47073
rect 3973 47107 4031 47113
rect 3973 47073 3985 47107
rect 4019 47104 4031 47107
rect 4890 47104 4896 47116
rect 4019 47076 4896 47104
rect 4019 47073 4031 47076
rect 3973 47067 4031 47073
rect 4890 47064 4896 47076
rect 4948 47064 4954 47116
rect 5166 47104 5172 47116
rect 5127 47076 5172 47104
rect 5166 47064 5172 47076
rect 5224 47064 5230 47116
rect 6564 47113 6592 47144
rect 20806 47132 20812 47184
rect 20864 47172 20870 47184
rect 20901 47175 20959 47181
rect 20901 47172 20913 47175
rect 20864 47144 20913 47172
rect 20864 47132 20870 47144
rect 20901 47141 20913 47144
rect 20947 47141 20959 47175
rect 20901 47135 20959 47141
rect 6549 47107 6607 47113
rect 6549 47073 6561 47107
rect 6595 47073 6607 47107
rect 6549 47067 6607 47073
rect 7374 47064 7380 47116
rect 7432 47104 7438 47116
rect 8389 47107 8447 47113
rect 8389 47104 8401 47107
rect 7432 47076 8401 47104
rect 7432 47064 7438 47076
rect 8389 47073 8401 47076
rect 8435 47073 8447 47107
rect 17402 47104 17408 47116
rect 17363 47076 17408 47104
rect 8389 47067 8447 47073
rect 17402 47064 17408 47076
rect 17460 47064 17466 47116
rect 29730 47064 29736 47116
rect 29788 47104 29794 47116
rect 30009 47107 30067 47113
rect 30009 47104 30021 47107
rect 29788 47076 30021 47104
rect 29788 47064 29794 47076
rect 30009 47073 30021 47076
rect 30055 47073 30067 47107
rect 30009 47067 30067 47073
rect 32306 47064 32312 47116
rect 32364 47104 32370 47116
rect 32585 47107 32643 47113
rect 32585 47104 32597 47107
rect 32364 47076 32597 47104
rect 32364 47064 32370 47076
rect 32585 47073 32597 47076
rect 32631 47073 32643 47107
rect 32585 47067 32643 47073
rect 35989 47107 36047 47113
rect 35989 47073 36001 47107
rect 36035 47104 36047 47107
rect 36722 47104 36728 47116
rect 36035 47076 36728 47104
rect 36035 47073 36047 47076
rect 35989 47067 36047 47073
rect 36722 47064 36728 47076
rect 36780 47064 36786 47116
rect 8938 47036 8944 47048
rect 8899 47008 8944 47036
rect 8938 46996 8944 47008
rect 8996 46996 9002 47048
rect 9766 47036 9772 47048
rect 9727 47008 9772 47036
rect 9766 46996 9772 47008
rect 9824 46996 9830 47048
rect 16850 47036 16856 47048
rect 16811 47008 16856 47036
rect 16850 46996 16856 47008
rect 16908 46996 16914 47048
rect 20162 46996 20168 47048
rect 20220 47036 20226 47048
rect 20257 47039 20315 47045
rect 20257 47036 20269 47039
rect 20220 47008 20269 47036
rect 20220 46996 20226 47008
rect 20257 47005 20269 47008
rect 20303 47005 20315 47039
rect 21085 47039 21143 47045
rect 21085 47036 21097 47039
rect 20257 46999 20315 47005
rect 20732 47008 21097 47036
rect 3050 46968 3056 46980
rect 3011 46940 3056 46968
rect 3050 46928 3056 46940
rect 3108 46928 3114 46980
rect 4157 46971 4215 46977
rect 4157 46937 4169 46971
rect 4203 46968 4215 46971
rect 4614 46968 4620 46980
rect 4203 46940 4620 46968
rect 4203 46937 4215 46940
rect 4157 46931 4215 46937
rect 4614 46928 4620 46940
rect 4672 46928 4678 46980
rect 8202 46968 8208 46980
rect 8163 46940 8208 46968
rect 8202 46928 8208 46940
rect 8260 46928 8266 46980
rect 17034 46968 17040 46980
rect 16995 46940 17040 46968
rect 17034 46928 17040 46940
rect 17092 46928 17098 46980
rect 19978 46860 19984 46912
rect 20036 46900 20042 46912
rect 20732 46900 20760 47008
rect 21085 47005 21097 47008
rect 21131 47005 21143 47039
rect 21085 46999 21143 47005
rect 22094 46996 22100 47048
rect 22152 47036 22158 47048
rect 22189 47039 22247 47045
rect 22189 47036 22201 47039
rect 22152 47008 22201 47036
rect 22152 46996 22158 47008
rect 22189 47005 22201 47008
rect 22235 47005 22247 47039
rect 24394 47036 24400 47048
rect 24355 47008 24400 47036
rect 22189 46999 22247 47005
rect 24394 46996 24400 47008
rect 24452 46996 24458 47048
rect 27982 47036 27988 47048
rect 27943 47008 27988 47036
rect 27982 46996 27988 47008
rect 28040 46996 28046 47048
rect 29546 47036 29552 47048
rect 29507 47008 29552 47036
rect 29546 46996 29552 47008
rect 29604 46996 29610 47048
rect 32122 47036 32128 47048
rect 32083 47008 32128 47036
rect 32122 46996 32128 47008
rect 32180 46996 32186 47048
rect 36446 47036 36452 47048
rect 36407 47008 36452 47036
rect 36446 46996 36452 47008
rect 36504 46996 36510 47048
rect 37734 47036 37740 47048
rect 37695 47008 37740 47036
rect 37734 46996 37740 47008
rect 37792 46996 37798 47048
rect 29270 46928 29276 46980
rect 29328 46968 29334 46980
rect 29733 46971 29791 46977
rect 29733 46968 29745 46971
rect 29328 46940 29745 46968
rect 29328 46928 29334 46940
rect 29733 46937 29745 46940
rect 29779 46937 29791 46971
rect 32306 46968 32312 46980
rect 32267 46940 32312 46968
rect 29733 46931 29791 46937
rect 32306 46928 32312 46940
rect 32364 46928 32370 46980
rect 20036 46872 20760 46900
rect 20036 46860 20042 46872
rect 1104 46810 38824 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 38824 46810
rect 1104 46736 38824 46758
rect 7377 46699 7435 46705
rect 7377 46665 7389 46699
rect 7423 46696 7435 46699
rect 8202 46696 8208 46708
rect 7423 46668 8208 46696
rect 7423 46665 7435 46668
rect 7377 46659 7435 46665
rect 8202 46656 8208 46668
rect 8260 46656 8266 46708
rect 2590 46588 2596 46640
rect 2648 46628 2654 46640
rect 7929 46631 7987 46637
rect 2648 46600 4384 46628
rect 2648 46588 2654 46600
rect 4356 46569 4384 46600
rect 7929 46597 7941 46631
rect 7975 46628 7987 46631
rect 8386 46628 8392 46640
rect 7975 46600 8392 46628
rect 7975 46597 7987 46600
rect 7929 46591 7987 46597
rect 8386 46588 8392 46600
rect 8444 46588 8450 46640
rect 33226 46628 33232 46640
rect 20548 46600 33232 46628
rect 20548 46572 20576 46600
rect 33226 46588 33232 46600
rect 33284 46588 33290 46640
rect 34425 46631 34483 46637
rect 34425 46597 34437 46631
rect 34471 46628 34483 46631
rect 35342 46628 35348 46640
rect 34471 46600 35348 46628
rect 34471 46597 34483 46600
rect 34425 46591 34483 46597
rect 35342 46588 35348 46600
rect 35400 46588 35406 46640
rect 36541 46631 36599 46637
rect 36541 46597 36553 46631
rect 36587 46628 36599 46631
rect 37553 46631 37611 46637
rect 37553 46628 37565 46631
rect 36587 46600 37565 46628
rect 36587 46597 36599 46600
rect 36541 46591 36599 46597
rect 37553 46597 37565 46600
rect 37599 46597 37611 46631
rect 37553 46591 37611 46597
rect 4341 46563 4399 46569
rect 4341 46529 4353 46563
rect 4387 46529 4399 46563
rect 4341 46523 4399 46529
rect 7469 46563 7527 46569
rect 7469 46529 7481 46563
rect 7515 46560 7527 46563
rect 8110 46560 8116 46572
rect 7515 46532 8116 46560
rect 7515 46529 7527 46532
rect 7469 46523 7527 46529
rect 8110 46520 8116 46532
rect 8168 46520 8174 46572
rect 9766 46520 9772 46572
rect 9824 46560 9830 46572
rect 9824 46532 9869 46560
rect 9824 46520 9830 46532
rect 16850 46520 16856 46572
rect 16908 46560 16914 46572
rect 16945 46563 17003 46569
rect 16945 46560 16957 46563
rect 16908 46532 16957 46560
rect 16908 46520 16914 46532
rect 16945 46529 16957 46532
rect 16991 46529 17003 46563
rect 20530 46560 20536 46572
rect 20491 46532 20536 46560
rect 16945 46523 17003 46529
rect 20530 46520 20536 46532
rect 20588 46520 20594 46572
rect 21174 46560 21180 46572
rect 21135 46532 21180 46560
rect 21174 46520 21180 46532
rect 21232 46520 21238 46572
rect 22094 46560 22100 46572
rect 22055 46532 22100 46560
rect 22094 46520 22100 46532
rect 22152 46520 22158 46572
rect 24394 46560 24400 46572
rect 24355 46532 24400 46560
rect 24394 46520 24400 46532
rect 24452 46520 24458 46572
rect 27982 46560 27988 46572
rect 27943 46532 27988 46560
rect 27982 46520 27988 46532
rect 28040 46520 28046 46572
rect 30469 46563 30527 46569
rect 30469 46529 30481 46563
rect 30515 46560 30527 46563
rect 32122 46560 32128 46572
rect 30515 46532 32128 46560
rect 30515 46529 30527 46532
rect 30469 46523 30527 46529
rect 32122 46520 32128 46532
rect 32180 46520 32186 46572
rect 36722 46520 36728 46572
rect 36780 46560 36786 46572
rect 37461 46563 37519 46569
rect 36780 46532 36825 46560
rect 36780 46520 36786 46532
rect 37461 46529 37473 46563
rect 37507 46560 37519 46563
rect 38010 46560 38016 46572
rect 37507 46532 38016 46560
rect 37507 46529 37519 46532
rect 37461 46523 37519 46529
rect 38010 46520 38016 46532
rect 38068 46520 38074 46572
rect 1581 46495 1639 46501
rect 1581 46461 1593 46495
rect 1627 46492 1639 46495
rect 2041 46495 2099 46501
rect 2041 46492 2053 46495
rect 1627 46464 2053 46492
rect 1627 46461 1639 46464
rect 1581 46455 1639 46461
rect 2041 46461 2053 46464
rect 2087 46461 2099 46495
rect 2041 46455 2099 46461
rect 2225 46495 2283 46501
rect 2225 46461 2237 46495
rect 2271 46492 2283 46495
rect 2774 46492 2780 46504
rect 2271 46464 2780 46492
rect 2271 46461 2283 46464
rect 2225 46455 2283 46461
rect 2774 46452 2780 46464
rect 2832 46452 2838 46504
rect 2958 46492 2964 46504
rect 2919 46464 2964 46492
rect 2958 46452 2964 46464
rect 3016 46452 3022 46504
rect 4617 46495 4675 46501
rect 4617 46461 4629 46495
rect 4663 46492 4675 46495
rect 5442 46492 5448 46504
rect 4663 46464 5448 46492
rect 4663 46461 4675 46464
rect 4617 46455 4675 46461
rect 5442 46452 5448 46464
rect 5500 46452 5506 46504
rect 8202 46452 8208 46504
rect 8260 46492 8266 46504
rect 9585 46495 9643 46501
rect 9585 46492 9597 46495
rect 8260 46464 9597 46492
rect 8260 46452 8266 46464
rect 9585 46461 9597 46464
rect 9631 46461 9643 46495
rect 9585 46455 9643 46461
rect 17589 46495 17647 46501
rect 17589 46461 17601 46495
rect 17635 46492 17647 46495
rect 18049 46495 18107 46501
rect 18049 46492 18061 46495
rect 17635 46464 18061 46492
rect 17635 46461 17647 46464
rect 17589 46455 17647 46461
rect 18049 46461 18061 46464
rect 18095 46461 18107 46495
rect 18230 46492 18236 46504
rect 18191 46464 18236 46492
rect 18049 46455 18107 46461
rect 18230 46452 18236 46464
rect 18288 46452 18294 46504
rect 18690 46492 18696 46504
rect 18651 46464 18696 46492
rect 18690 46452 18696 46464
rect 18748 46452 18754 46504
rect 22281 46495 22339 46501
rect 22281 46461 22293 46495
rect 22327 46492 22339 46495
rect 22554 46492 22560 46504
rect 22327 46464 22560 46492
rect 22327 46461 22339 46464
rect 22281 46455 22339 46461
rect 22554 46452 22560 46464
rect 22612 46452 22618 46504
rect 22646 46452 22652 46504
rect 22704 46492 22710 46504
rect 24578 46492 24584 46504
rect 22704 46464 22749 46492
rect 24539 46464 24584 46492
rect 22704 46452 22710 46464
rect 24578 46452 24584 46464
rect 24636 46452 24642 46504
rect 24857 46495 24915 46501
rect 24857 46461 24869 46495
rect 24903 46461 24915 46495
rect 24857 46455 24915 46461
rect 28169 46495 28227 46501
rect 28169 46461 28181 46495
rect 28215 46492 28227 46495
rect 28626 46492 28632 46504
rect 28215 46464 28632 46492
rect 28215 46461 28227 46464
rect 28169 46455 28227 46461
rect 24486 46384 24492 46436
rect 24544 46424 24550 46436
rect 24872 46424 24900 46455
rect 28626 46452 28632 46464
rect 28684 46452 28690 46504
rect 28721 46495 28779 46501
rect 28721 46461 28733 46495
rect 28767 46461 28779 46495
rect 28721 46455 28779 46461
rect 32585 46495 32643 46501
rect 32585 46461 32597 46495
rect 32631 46461 32643 46495
rect 32585 46455 32643 46461
rect 32769 46495 32827 46501
rect 32769 46461 32781 46495
rect 32815 46492 32827 46495
rect 33318 46492 33324 46504
rect 32815 46464 33324 46492
rect 32815 46461 32827 46464
rect 32769 46455 32827 46461
rect 24544 46396 24900 46424
rect 24544 46384 24550 46396
rect 28350 46384 28356 46436
rect 28408 46424 28414 46436
rect 28736 46424 28764 46455
rect 28408 46396 28764 46424
rect 32600 46424 32628 46455
rect 33318 46452 33324 46464
rect 33376 46452 33382 46504
rect 35802 46492 35808 46504
rect 35763 46464 35808 46492
rect 35802 46452 35808 46464
rect 35860 46452 35866 46504
rect 33870 46424 33876 46436
rect 32600 46396 33876 46424
rect 28408 46384 28414 46396
rect 33870 46384 33876 46396
rect 33928 46384 33934 46436
rect 5810 46356 5816 46368
rect 5771 46328 5816 46356
rect 5810 46316 5816 46328
rect 5868 46316 5874 46368
rect 6086 46316 6092 46368
rect 6144 46356 6150 46368
rect 6365 46359 6423 46365
rect 6365 46356 6377 46359
rect 6144 46328 6377 46356
rect 6144 46316 6150 46328
rect 6365 46325 6377 46328
rect 6411 46325 6423 46359
rect 6365 46319 6423 46325
rect 14918 46316 14924 46368
rect 14976 46356 14982 46368
rect 15013 46359 15071 46365
rect 15013 46356 15025 46359
rect 14976 46328 15025 46356
rect 14976 46316 14982 46328
rect 15013 46325 15025 46328
rect 15059 46325 15071 46359
rect 15013 46319 15071 46325
rect 16117 46359 16175 46365
rect 16117 46325 16129 46359
rect 16163 46356 16175 46359
rect 19426 46356 19432 46368
rect 16163 46328 19432 46356
rect 16163 46325 16175 46328
rect 16117 46319 16175 46325
rect 19426 46316 19432 46328
rect 19484 46316 19490 46368
rect 20346 46316 20352 46368
rect 20404 46356 20410 46368
rect 20441 46359 20499 46365
rect 20441 46356 20453 46359
rect 20404 46328 20453 46356
rect 20404 46316 20410 46328
rect 20441 46325 20453 46328
rect 20487 46325 20499 46359
rect 20441 46319 20499 46325
rect 20993 46359 21051 46365
rect 20993 46325 21005 46359
rect 21039 46356 21051 46359
rect 21082 46356 21088 46368
rect 21039 46328 21088 46356
rect 21039 46325 21051 46328
rect 20993 46319 21051 46325
rect 21082 46316 21088 46328
rect 21140 46316 21146 46368
rect 26234 46316 26240 46368
rect 26292 46356 26298 46368
rect 26973 46359 27031 46365
rect 26973 46356 26985 46359
rect 26292 46328 26985 46356
rect 26292 46316 26298 46328
rect 26973 46325 26985 46328
rect 27019 46325 27031 46359
rect 30926 46356 30932 46368
rect 30887 46328 30932 46356
rect 26973 46319 27031 46325
rect 30926 46316 30932 46328
rect 30984 46316 30990 46368
rect 1104 46266 38824 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 38824 46266
rect 1104 46192 38824 46214
rect 3050 46112 3056 46164
rect 3108 46152 3114 46164
rect 3881 46155 3939 46161
rect 3881 46152 3893 46155
rect 3108 46124 3893 46152
rect 3108 46112 3114 46124
rect 3881 46121 3893 46124
rect 3927 46121 3939 46155
rect 4614 46152 4620 46164
rect 4575 46124 4620 46152
rect 3881 46115 3939 46121
rect 4614 46112 4620 46124
rect 4672 46112 4678 46164
rect 4890 46112 4896 46164
rect 4948 46152 4954 46164
rect 5169 46155 5227 46161
rect 5169 46152 5181 46155
rect 4948 46124 5181 46152
rect 4948 46112 4954 46124
rect 5169 46121 5181 46124
rect 5215 46121 5227 46155
rect 8202 46152 8208 46164
rect 8163 46124 8208 46152
rect 5169 46115 5227 46121
rect 8202 46112 8208 46124
rect 8260 46112 8266 46164
rect 17034 46112 17040 46164
rect 17092 46152 17098 46164
rect 17313 46155 17371 46161
rect 17313 46152 17325 46155
rect 17092 46124 17325 46152
rect 17092 46112 17098 46124
rect 17313 46121 17325 46124
rect 17359 46121 17371 46155
rect 18230 46152 18236 46164
rect 18191 46124 18236 46152
rect 17313 46115 17371 46121
rect 18230 46112 18236 46124
rect 18288 46112 18294 46164
rect 22554 46152 22560 46164
rect 22515 46124 22560 46152
rect 22554 46112 22560 46124
rect 22612 46112 22618 46164
rect 24489 46155 24547 46161
rect 24489 46121 24501 46155
rect 24535 46152 24547 46155
rect 24578 46152 24584 46164
rect 24535 46124 24584 46152
rect 24535 46121 24547 46124
rect 24489 46115 24547 46121
rect 24578 46112 24584 46124
rect 24636 46112 24642 46164
rect 28626 46152 28632 46164
rect 28587 46124 28632 46152
rect 28626 46112 28632 46124
rect 28684 46112 28690 46164
rect 29546 46152 29552 46164
rect 29507 46124 29552 46152
rect 29546 46112 29552 46124
rect 29604 46112 29610 46164
rect 33318 46152 33324 46164
rect 33279 46124 33324 46152
rect 33318 46112 33324 46124
rect 33376 46112 33382 46164
rect 33870 46152 33876 46164
rect 33831 46124 33876 46152
rect 33870 46112 33876 46124
rect 33928 46112 33934 46164
rect 9030 46044 9036 46096
rect 9088 46044 9094 46096
rect 14 45976 20 46028
rect 72 46016 78 46028
rect 1397 46019 1455 46025
rect 1397 46016 1409 46019
rect 72 45988 1409 46016
rect 72 45976 78 45988
rect 1397 45985 1409 45988
rect 1443 45985 1455 46019
rect 1397 45979 1455 45985
rect 5813 46019 5871 46025
rect 5813 45985 5825 46019
rect 5859 46016 5871 46019
rect 6086 46016 6092 46028
rect 5859 45988 6092 46016
rect 5859 45985 5871 45988
rect 5813 45979 5871 45985
rect 6086 45976 6092 45988
rect 6144 45976 6150 46028
rect 6454 46016 6460 46028
rect 6415 45988 6460 46016
rect 6454 45976 6460 45988
rect 6512 45976 6518 46028
rect 8938 46016 8944 46028
rect 8899 45988 8944 46016
rect 8938 45976 8944 45988
rect 8996 45976 9002 46028
rect 9048 46016 9076 46044
rect 9401 46019 9459 46025
rect 9401 46016 9413 46019
rect 9048 45988 9413 46016
rect 9401 45985 9413 45988
rect 9447 45985 9459 46019
rect 14918 46016 14924 46028
rect 14879 45988 14924 46016
rect 9401 45979 9459 45985
rect 14918 45976 14924 45988
rect 14976 45976 14982 46028
rect 15470 46016 15476 46028
rect 15431 45988 15476 46016
rect 15470 45976 15476 45988
rect 15528 45976 15534 46028
rect 20162 46016 20168 46028
rect 17420 45988 19472 46016
rect 20123 45988 20168 46016
rect 17420 45960 17448 45988
rect 3234 45908 3240 45960
rect 3292 45948 3298 45960
rect 3973 45951 4031 45957
rect 3292 45920 3337 45948
rect 3292 45908 3298 45920
rect 3973 45917 3985 45951
rect 4019 45948 4031 45951
rect 4709 45951 4767 45957
rect 4709 45948 4721 45951
rect 4019 45920 4721 45948
rect 4019 45917 4031 45920
rect 3973 45911 4031 45917
rect 4709 45917 4721 45920
rect 4755 45948 4767 45951
rect 4798 45948 4804 45960
rect 4755 45920 4804 45948
rect 4755 45917 4767 45920
rect 4709 45911 4767 45917
rect 4798 45908 4804 45920
rect 4856 45908 4862 45960
rect 8110 45948 8116 45960
rect 8071 45920 8116 45948
rect 8110 45908 8116 45920
rect 8168 45908 8174 45960
rect 17402 45948 17408 45960
rect 17363 45920 17408 45948
rect 17402 45908 17408 45920
rect 17460 45908 17466 45960
rect 18046 45908 18052 45960
rect 18104 45948 18110 45960
rect 19444 45957 19472 45988
rect 20162 45976 20168 45988
rect 20220 45976 20226 46028
rect 20346 46016 20352 46028
rect 20307 45988 20352 46016
rect 20346 45976 20352 45988
rect 20404 45976 20410 46028
rect 21266 46016 21272 46028
rect 21227 45988 21272 46016
rect 21266 45976 21272 45988
rect 21324 45976 21330 46028
rect 26234 45976 26240 46028
rect 26292 46016 26298 46028
rect 27062 46016 27068 46028
rect 26292 45988 26337 46016
rect 27023 45988 27068 46016
rect 26292 45976 26298 45988
rect 27062 45976 27068 45988
rect 27120 45976 27126 46028
rect 30926 46016 30932 46028
rect 30887 45988 30932 46016
rect 30926 45976 30932 45988
rect 30984 45976 30990 46028
rect 31570 45976 31576 46028
rect 31628 46016 31634 46028
rect 31757 46019 31815 46025
rect 31757 46016 31769 46019
rect 31628 45988 31769 46016
rect 31628 45976 31634 45988
rect 31757 45985 31769 45988
rect 31803 45985 31815 46019
rect 31757 45979 31815 45985
rect 36265 46019 36323 46025
rect 36265 45985 36277 46019
rect 36311 46016 36323 46019
rect 36446 46016 36452 46028
rect 36311 45988 36452 46016
rect 36311 45985 36323 45988
rect 36265 45979 36323 45985
rect 36446 45976 36452 45988
rect 36504 45976 36510 46028
rect 37366 46016 37372 46028
rect 37327 45988 37372 46016
rect 37366 45976 37372 45988
rect 37424 45976 37430 46028
rect 18141 45951 18199 45957
rect 18141 45948 18153 45951
rect 18104 45920 18153 45948
rect 18104 45908 18110 45920
rect 18141 45917 18153 45920
rect 18187 45917 18199 45951
rect 18141 45911 18199 45917
rect 19429 45951 19487 45957
rect 19429 45917 19441 45951
rect 19475 45917 19487 45951
rect 22646 45948 22652 45960
rect 22607 45920 22652 45948
rect 19429 45911 19487 45917
rect 22646 45908 22652 45920
rect 22704 45908 22710 45960
rect 23842 45908 23848 45960
rect 23900 45948 23906 45960
rect 24397 45951 24455 45957
rect 24397 45948 24409 45951
rect 23900 45920 24409 45948
rect 23900 45908 23906 45920
rect 24397 45917 24409 45920
rect 24443 45948 24455 45951
rect 28718 45948 28724 45960
rect 24443 45920 26234 45948
rect 28679 45920 28724 45948
rect 24443 45917 24455 45920
rect 24397 45911 24455 45917
rect 3050 45880 3056 45892
rect 3011 45852 3056 45880
rect 3050 45840 3056 45852
rect 3108 45840 3114 45892
rect 5718 45840 5724 45892
rect 5776 45880 5782 45892
rect 5997 45883 6055 45889
rect 5997 45880 6009 45883
rect 5776 45852 6009 45880
rect 5776 45840 5782 45852
rect 5997 45849 6009 45852
rect 6043 45849 6055 45883
rect 5997 45843 6055 45849
rect 8938 45840 8944 45892
rect 8996 45880 9002 45892
rect 9125 45883 9183 45889
rect 9125 45880 9137 45883
rect 8996 45852 9137 45880
rect 8996 45840 9002 45852
rect 9125 45849 9137 45852
rect 9171 45849 9183 45883
rect 9125 45843 9183 45849
rect 15105 45883 15163 45889
rect 15105 45849 15117 45883
rect 15151 45880 15163 45883
rect 15194 45880 15200 45892
rect 15151 45852 15200 45880
rect 15151 45849 15163 45852
rect 15105 45843 15163 45849
rect 15194 45840 15200 45852
rect 15252 45840 15258 45892
rect 7466 45772 7472 45824
rect 7524 45812 7530 45824
rect 8110 45812 8116 45824
rect 7524 45784 8116 45812
rect 7524 45772 7530 45784
rect 8110 45772 8116 45784
rect 8168 45772 8174 45824
rect 19334 45812 19340 45824
rect 19295 45784 19340 45812
rect 19334 45772 19340 45784
rect 19392 45772 19398 45824
rect 26206 45812 26234 45920
rect 28718 45908 28724 45920
rect 28776 45908 28782 45960
rect 33226 45948 33232 45960
rect 33187 45920 33232 45948
rect 33226 45908 33232 45920
rect 33284 45908 33290 45960
rect 26418 45880 26424 45892
rect 26379 45852 26424 45880
rect 26418 45840 26424 45852
rect 26476 45840 26482 45892
rect 31110 45880 31116 45892
rect 31071 45852 31116 45880
rect 31110 45840 31116 45852
rect 31168 45840 31174 45892
rect 36449 45883 36507 45889
rect 36449 45849 36461 45883
rect 36495 45880 36507 45883
rect 37366 45880 37372 45892
rect 36495 45852 37372 45880
rect 36495 45849 36507 45852
rect 36449 45843 36507 45849
rect 37366 45840 37372 45852
rect 37424 45840 37430 45892
rect 38010 45812 38016 45824
rect 26206 45784 38016 45812
rect 38010 45772 38016 45784
rect 38068 45772 38074 45824
rect 1104 45722 38824 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 38824 45722
rect 1104 45648 38824 45670
rect 5718 45608 5724 45620
rect 5679 45580 5724 45608
rect 5718 45568 5724 45580
rect 5776 45568 5782 45620
rect 8938 45608 8944 45620
rect 8899 45580 8944 45608
rect 8938 45568 8944 45580
rect 8996 45568 9002 45620
rect 25317 45611 25375 45617
rect 25317 45577 25329 45611
rect 25363 45608 25375 45611
rect 26329 45611 26387 45617
rect 25363 45580 25397 45608
rect 25363 45577 25375 45580
rect 25317 45571 25375 45577
rect 26329 45577 26341 45611
rect 26375 45608 26387 45611
rect 26418 45608 26424 45620
rect 26375 45580 26424 45608
rect 26375 45577 26387 45580
rect 26329 45571 26387 45577
rect 2774 45540 2780 45552
rect 2735 45512 2780 45540
rect 2774 45500 2780 45512
rect 2832 45500 2838 45552
rect 6914 45540 6920 45552
rect 5644 45512 6920 45540
rect 2869 45475 2927 45481
rect 2869 45441 2881 45475
rect 2915 45472 2927 45475
rect 2958 45472 2964 45484
rect 2915 45444 2964 45472
rect 2915 45441 2927 45444
rect 2869 45435 2927 45441
rect 2958 45432 2964 45444
rect 3016 45432 3022 45484
rect 3234 45432 3240 45484
rect 3292 45472 3298 45484
rect 5644 45481 5672 45512
rect 6914 45500 6920 45512
rect 6972 45500 6978 45552
rect 15194 45540 15200 45552
rect 15155 45512 15200 45540
rect 15194 45500 15200 45512
rect 15252 45500 15258 45552
rect 19153 45543 19211 45549
rect 19153 45509 19165 45543
rect 19199 45540 19211 45543
rect 19334 45540 19340 45552
rect 19199 45512 19340 45540
rect 19199 45509 19211 45512
rect 19153 45503 19211 45509
rect 19334 45500 19340 45512
rect 19392 45500 19398 45552
rect 24612 45543 24670 45549
rect 20824 45512 23612 45540
rect 3329 45475 3387 45481
rect 3329 45472 3341 45475
rect 3292 45444 3341 45472
rect 3292 45432 3298 45444
rect 3329 45441 3341 45444
rect 3375 45441 3387 45475
rect 3329 45435 3387 45441
rect 5629 45475 5687 45481
rect 5629 45441 5641 45475
rect 5675 45441 5687 45475
rect 5629 45435 5687 45441
rect 5810 45432 5816 45484
rect 5868 45472 5874 45484
rect 6549 45475 6607 45481
rect 6549 45472 6561 45475
rect 5868 45444 6561 45472
rect 5868 45432 5874 45444
rect 6549 45441 6561 45444
rect 6595 45441 6607 45475
rect 6549 45435 6607 45441
rect 8018 45432 8024 45484
rect 8076 45472 8082 45484
rect 8076 45444 8800 45472
rect 8076 45432 8082 45444
rect 1394 45404 1400 45416
rect 1355 45376 1400 45404
rect 1394 45364 1400 45376
rect 1452 45364 1458 45416
rect 1670 45404 1676 45416
rect 1631 45376 1676 45404
rect 1670 45364 1676 45376
rect 1728 45364 1734 45416
rect 6730 45404 6736 45416
rect 6691 45376 6736 45404
rect 6730 45364 6736 45376
rect 6788 45364 6794 45416
rect 8110 45404 8116 45416
rect 8071 45376 8116 45404
rect 8110 45364 8116 45376
rect 8168 45364 8174 45416
rect 8772 45404 8800 45444
rect 8846 45432 8852 45484
rect 8904 45472 8910 45484
rect 15286 45472 15292 45484
rect 8904 45444 8949 45472
rect 15247 45444 15292 45472
rect 8904 45432 8910 45444
rect 15286 45432 15292 45444
rect 15344 45432 15350 45484
rect 20070 45481 20076 45484
rect 20064 45435 20076 45481
rect 20128 45472 20134 45484
rect 20128 45444 20164 45472
rect 20070 45432 20076 45435
rect 20128 45432 20134 45444
rect 17954 45404 17960 45416
rect 8772 45376 12434 45404
rect 17915 45376 17960 45404
rect 2958 45296 2964 45348
rect 3016 45336 3022 45348
rect 10042 45336 10048 45348
rect 3016 45308 10048 45336
rect 3016 45296 3022 45308
rect 10042 45296 10048 45308
rect 10100 45296 10106 45348
rect 12406 45268 12434 45376
rect 17954 45364 17960 45376
rect 18012 45364 18018 45416
rect 19337 45407 19395 45413
rect 19337 45373 19349 45407
rect 19383 45404 19395 45407
rect 19426 45404 19432 45416
rect 19383 45376 19432 45404
rect 19383 45373 19395 45376
rect 19337 45367 19395 45373
rect 19426 45364 19432 45376
rect 19484 45364 19490 45416
rect 19794 45404 19800 45416
rect 19755 45376 19800 45404
rect 19794 45364 19800 45376
rect 19852 45364 19858 45416
rect 20824 45268 20852 45512
rect 22094 45432 22100 45484
rect 22152 45472 22158 45484
rect 22373 45475 22431 45481
rect 22373 45472 22385 45475
rect 22152 45444 22385 45472
rect 22152 45432 22158 45444
rect 22373 45441 22385 45444
rect 22419 45441 22431 45475
rect 22373 45435 22431 45441
rect 22649 45475 22707 45481
rect 22649 45441 22661 45475
rect 22695 45472 22707 45475
rect 23014 45472 23020 45484
rect 22695 45444 23020 45472
rect 22695 45441 22707 45444
rect 22649 45435 22707 45441
rect 23014 45432 23020 45444
rect 23072 45432 23078 45484
rect 22557 45407 22615 45413
rect 22557 45373 22569 45407
rect 22603 45373 22615 45407
rect 22557 45367 22615 45373
rect 22572 45336 22600 45367
rect 22922 45336 22928 45348
rect 22066 45308 22416 45336
rect 22572 45308 22928 45336
rect 12406 45240 20852 45268
rect 20898 45228 20904 45280
rect 20956 45268 20962 45280
rect 21177 45271 21235 45277
rect 21177 45268 21189 45271
rect 20956 45240 21189 45268
rect 20956 45228 20962 45240
rect 21177 45237 21189 45240
rect 21223 45268 21235 45271
rect 22066 45268 22094 45308
rect 22186 45268 22192 45280
rect 21223 45240 22094 45268
rect 22147 45240 22192 45268
rect 21223 45237 21235 45240
rect 21177 45231 21235 45237
rect 22186 45228 22192 45240
rect 22244 45228 22250 45280
rect 22388 45277 22416 45308
rect 22922 45296 22928 45308
rect 22980 45336 22986 45348
rect 23477 45339 23535 45345
rect 23477 45336 23489 45339
rect 22980 45308 23489 45336
rect 22980 45296 22986 45308
rect 23477 45305 23489 45308
rect 23523 45305 23535 45339
rect 23477 45299 23535 45305
rect 22373 45271 22431 45277
rect 22373 45237 22385 45271
rect 22419 45268 22431 45271
rect 22830 45268 22836 45280
rect 22419 45240 22836 45268
rect 22419 45237 22431 45240
rect 22373 45231 22431 45237
rect 22830 45228 22836 45240
rect 22888 45228 22894 45280
rect 23584 45268 23612 45512
rect 24612 45509 24624 45543
rect 24658 45540 24670 45543
rect 25332 45540 25360 45571
rect 26418 45568 26424 45580
rect 26476 45568 26482 45620
rect 31110 45608 31116 45620
rect 31071 45580 31116 45608
rect 31110 45568 31116 45580
rect 31168 45568 31174 45620
rect 29270 45540 29276 45552
rect 24658 45512 25360 45540
rect 29231 45512 29276 45540
rect 24658 45509 24670 45512
rect 24612 45503 24670 45509
rect 29270 45500 29276 45512
rect 29328 45500 29334 45552
rect 32217 45543 32275 45549
rect 32217 45509 32229 45543
rect 32263 45540 32275 45543
rect 32306 45540 32312 45552
rect 32263 45512 32312 45540
rect 32263 45509 32275 45512
rect 32217 45503 32275 45509
rect 32306 45500 32312 45512
rect 32364 45500 32370 45552
rect 37366 45540 37372 45552
rect 37327 45512 37372 45540
rect 37366 45500 37372 45512
rect 37424 45500 37430 45552
rect 24762 45432 24768 45484
rect 24820 45472 24826 45484
rect 24857 45475 24915 45481
rect 24857 45472 24869 45475
rect 24820 45444 24869 45472
rect 24820 45432 24826 45444
rect 24857 45441 24869 45444
rect 24903 45441 24915 45475
rect 24857 45435 24915 45441
rect 24946 45432 24952 45484
rect 25004 45472 25010 45484
rect 25501 45475 25559 45481
rect 25501 45472 25513 45475
rect 25004 45444 25513 45472
rect 25004 45432 25010 45444
rect 25501 45441 25513 45444
rect 25547 45441 25559 45475
rect 25501 45435 25559 45441
rect 26237 45475 26295 45481
rect 26237 45441 26249 45475
rect 26283 45441 26295 45475
rect 26237 45435 26295 45441
rect 26252 45268 26280 45435
rect 27154 45432 27160 45484
rect 27212 45472 27218 45484
rect 28086 45475 28144 45481
rect 28086 45472 28098 45475
rect 27212 45444 28098 45472
rect 27212 45432 27218 45444
rect 28086 45441 28098 45444
rect 28132 45441 28144 45475
rect 28086 45435 28144 45441
rect 29181 45475 29239 45481
rect 29181 45441 29193 45475
rect 29227 45472 29239 45475
rect 31021 45475 31079 45481
rect 29227 45444 29316 45472
rect 29227 45441 29239 45444
rect 29181 45435 29239 45441
rect 29288 45416 29316 45444
rect 31021 45441 31033 45475
rect 31067 45472 31079 45475
rect 31202 45472 31208 45484
rect 31067 45444 31208 45472
rect 31067 45441 31079 45444
rect 31021 45435 31079 45441
rect 31202 45432 31208 45444
rect 31260 45432 31266 45484
rect 32125 45475 32183 45481
rect 32125 45441 32137 45475
rect 32171 45472 32183 45475
rect 32398 45472 32404 45484
rect 32171 45444 32404 45472
rect 32171 45441 32183 45444
rect 32125 45435 32183 45441
rect 32398 45432 32404 45444
rect 32456 45432 32462 45484
rect 37274 45472 37280 45484
rect 37235 45444 37280 45472
rect 37274 45432 37280 45444
rect 37332 45432 37338 45484
rect 37921 45475 37979 45481
rect 37921 45441 37933 45475
rect 37967 45472 37979 45475
rect 38378 45472 38384 45484
rect 37967 45444 38384 45472
rect 37967 45441 37979 45444
rect 37921 45435 37979 45441
rect 38378 45432 38384 45444
rect 38436 45432 38442 45484
rect 28350 45404 28356 45416
rect 28311 45376 28356 45404
rect 28350 45364 28356 45376
rect 28408 45364 28414 45416
rect 29270 45364 29276 45416
rect 29328 45364 29334 45416
rect 35802 45404 35808 45416
rect 35763 45376 35808 45404
rect 35802 45364 35808 45376
rect 35860 45364 35866 45416
rect 36538 45404 36544 45416
rect 36499 45376 36544 45404
rect 36538 45364 36544 45376
rect 36596 45364 36602 45416
rect 36722 45404 36728 45416
rect 36683 45376 36728 45404
rect 36722 45364 36728 45376
rect 36780 45364 36786 45416
rect 23584 45240 26280 45268
rect 26878 45228 26884 45280
rect 26936 45268 26942 45280
rect 26973 45271 27031 45277
rect 26973 45268 26985 45271
rect 26936 45240 26985 45268
rect 26936 45228 26942 45240
rect 26973 45237 26985 45240
rect 27019 45237 27031 45271
rect 26973 45231 27031 45237
rect 37918 45228 37924 45280
rect 37976 45268 37982 45280
rect 38013 45271 38071 45277
rect 38013 45268 38025 45271
rect 37976 45240 38025 45268
rect 37976 45228 37982 45240
rect 38013 45237 38025 45240
rect 38059 45237 38071 45271
rect 38013 45231 38071 45237
rect 1104 45178 38824 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 38824 45178
rect 1104 45104 38824 45126
rect 1765 45067 1823 45073
rect 1765 45033 1777 45067
rect 1811 45064 1823 45067
rect 2866 45064 2872 45076
rect 1811 45036 2872 45064
rect 1811 45033 1823 45036
rect 1765 45027 1823 45033
rect 2866 45024 2872 45036
rect 2924 45024 2930 45076
rect 6641 45067 6699 45073
rect 6641 45033 6653 45067
rect 6687 45064 6699 45067
rect 6730 45064 6736 45076
rect 6687 45036 6736 45064
rect 6687 45033 6699 45036
rect 6641 45027 6699 45033
rect 6730 45024 6736 45036
rect 6788 45024 6794 45076
rect 7374 45064 7380 45076
rect 7335 45036 7380 45064
rect 7374 45024 7380 45036
rect 7432 45024 7438 45076
rect 8846 45024 8852 45076
rect 8904 45064 8910 45076
rect 37366 45064 37372 45076
rect 8904 45036 37372 45064
rect 8904 45024 8910 45036
rect 37366 45024 37372 45036
rect 37424 45024 37430 45076
rect 2317 44999 2375 45005
rect 2317 44965 2329 44999
rect 2363 44996 2375 44999
rect 3050 44996 3056 45008
rect 2363 44968 3056 44996
rect 2363 44965 2375 44968
rect 2317 44959 2375 44965
rect 3050 44956 3056 44968
rect 3108 44956 3114 45008
rect 23014 44956 23020 45008
rect 23072 44996 23078 45008
rect 26697 44999 26755 45005
rect 23072 44968 24440 44996
rect 23072 44956 23078 44968
rect 18138 44888 18144 44940
rect 18196 44928 18202 44940
rect 19794 44928 19800 44940
rect 18196 44900 19800 44928
rect 18196 44888 18202 44900
rect 19794 44888 19800 44900
rect 19852 44928 19858 44940
rect 20809 44931 20867 44937
rect 20809 44928 20821 44931
rect 19852 44900 20821 44928
rect 19852 44888 19858 44900
rect 20809 44897 20821 44900
rect 20855 44897 20867 44931
rect 20809 44891 20867 44897
rect 2409 44863 2467 44869
rect 2409 44829 2421 44863
rect 2455 44860 2467 44863
rect 2498 44860 2504 44872
rect 2455 44832 2504 44860
rect 2455 44829 2467 44832
rect 2409 44823 2467 44829
rect 2498 44820 2504 44832
rect 2556 44820 2562 44872
rect 6549 44863 6607 44869
rect 6549 44829 6561 44863
rect 6595 44860 6607 44863
rect 6914 44860 6920 44872
rect 6595 44832 6920 44860
rect 6595 44829 6607 44832
rect 6549 44823 6607 44829
rect 6914 44820 6920 44832
rect 6972 44860 6978 44872
rect 8202 44860 8208 44872
rect 6972 44832 8208 44860
rect 6972 44820 6978 44832
rect 8202 44820 8208 44832
rect 8260 44820 8266 44872
rect 19426 44820 19432 44872
rect 19484 44860 19490 44872
rect 19521 44863 19579 44869
rect 19521 44860 19533 44863
rect 19484 44832 19533 44860
rect 19484 44820 19490 44832
rect 19521 44829 19533 44832
rect 19567 44829 19579 44863
rect 19521 44823 19579 44829
rect 19705 44863 19763 44869
rect 19705 44829 19717 44863
rect 19751 44860 19763 44863
rect 20714 44860 20720 44872
rect 19751 44832 20720 44860
rect 19751 44829 19763 44832
rect 19705 44823 19763 44829
rect 20714 44820 20720 44832
rect 20772 44820 20778 44872
rect 2498 44684 2504 44736
rect 2556 44724 2562 44736
rect 10502 44724 10508 44736
rect 2556 44696 10508 44724
rect 2556 44684 2562 44696
rect 10502 44684 10508 44696
rect 10560 44684 10566 44736
rect 19889 44727 19947 44733
rect 19889 44693 19901 44727
rect 19935 44724 19947 44727
rect 19978 44724 19984 44736
rect 19935 44696 19984 44724
rect 19935 44693 19947 44696
rect 19889 44687 19947 44693
rect 19978 44684 19984 44696
rect 20036 44684 20042 44736
rect 20824 44724 20852 44891
rect 22370 44888 22376 44940
rect 22428 44928 22434 44940
rect 24412 44937 24440 44968
rect 26697 44965 26709 44999
rect 26743 44996 26755 44999
rect 27338 44996 27344 45008
rect 26743 44968 27344 44996
rect 26743 44965 26755 44968
rect 26697 44959 26755 44965
rect 27338 44956 27344 44968
rect 27396 44996 27402 45008
rect 27396 44968 27568 44996
rect 27396 44956 27402 44968
rect 23201 44931 23259 44937
rect 23201 44928 23213 44931
rect 22428 44900 23213 44928
rect 22428 44888 22434 44900
rect 23201 44897 23213 44900
rect 23247 44897 23259 44931
rect 23201 44891 23259 44897
rect 24397 44931 24455 44937
rect 24397 44897 24409 44931
rect 24443 44897 24455 44931
rect 24397 44891 24455 44897
rect 24762 44888 24768 44940
rect 24820 44928 24826 44940
rect 27540 44937 27568 44968
rect 37734 44956 37740 45008
rect 37792 44996 37798 45008
rect 37792 44968 38148 44996
rect 37792 44956 37798 44968
rect 25317 44931 25375 44937
rect 25317 44928 25329 44931
rect 24820 44900 25329 44928
rect 24820 44888 24826 44900
rect 25317 44897 25329 44900
rect 25363 44897 25375 44931
rect 25317 44891 25375 44897
rect 27525 44931 27583 44937
rect 27525 44897 27537 44931
rect 27571 44897 27583 44931
rect 37090 44928 37096 44940
rect 37051 44900 37096 44928
rect 27525 44891 27583 44897
rect 37090 44888 37096 44900
rect 37148 44888 37154 44940
rect 37918 44928 37924 44940
rect 37879 44900 37924 44928
rect 37918 44888 37924 44900
rect 37976 44888 37982 44940
rect 38120 44937 38148 44968
rect 38105 44931 38163 44937
rect 38105 44897 38117 44931
rect 38151 44897 38163 44931
rect 38105 44891 38163 44897
rect 23566 44860 23572 44872
rect 21192 44832 23572 44860
rect 21082 44801 21088 44804
rect 21076 44792 21088 44801
rect 21043 44764 21088 44792
rect 21076 44755 21088 44764
rect 21082 44752 21088 44755
rect 21140 44752 21146 44804
rect 21192 44724 21220 44832
rect 23566 44820 23572 44832
rect 23624 44820 23630 44872
rect 23845 44863 23903 44869
rect 23845 44829 23857 44863
rect 23891 44829 23903 44863
rect 23845 44823 23903 44829
rect 24581 44863 24639 44869
rect 24581 44829 24593 44863
rect 24627 44860 24639 44863
rect 26050 44860 26056 44872
rect 24627 44832 26056 44860
rect 24627 44829 24639 44832
rect 24581 44823 24639 44829
rect 22649 44795 22707 44801
rect 22649 44761 22661 44795
rect 22695 44761 22707 44795
rect 22922 44792 22928 44804
rect 22883 44764 22928 44792
rect 22649 44755 22707 44761
rect 20824 44696 21220 44724
rect 22094 44684 22100 44736
rect 22152 44724 22158 44736
rect 22189 44727 22247 44733
rect 22189 44724 22201 44727
rect 22152 44696 22201 44724
rect 22152 44684 22158 44696
rect 22189 44693 22201 44696
rect 22235 44724 22247 44727
rect 22664 44724 22692 44755
rect 22922 44752 22928 44764
rect 22980 44752 22986 44804
rect 23106 44752 23112 44804
rect 23164 44792 23170 44804
rect 23860 44792 23888 44823
rect 26050 44820 26056 44832
rect 26108 44860 26114 44872
rect 27341 44863 27399 44869
rect 27341 44860 27353 44863
rect 26108 44832 27353 44860
rect 26108 44820 26114 44832
rect 27341 44829 27353 44832
rect 27387 44829 27399 44863
rect 27341 44823 27399 44829
rect 23164 44764 23888 44792
rect 24765 44795 24823 44801
rect 23164 44752 23170 44764
rect 24765 44761 24777 44795
rect 24811 44792 24823 44795
rect 24946 44792 24952 44804
rect 24811 44764 24952 44792
rect 24811 44761 24823 44764
rect 24765 44755 24823 44761
rect 24946 44752 24952 44764
rect 25004 44752 25010 44804
rect 25584 44795 25642 44801
rect 25584 44761 25596 44795
rect 25630 44792 25642 44795
rect 25774 44792 25780 44804
rect 25630 44764 25780 44792
rect 25630 44761 25642 44764
rect 25584 44755 25642 44761
rect 25774 44752 25780 44764
rect 25832 44752 25838 44804
rect 22830 44724 22836 44736
rect 22235 44696 22692 44724
rect 22791 44696 22836 44724
rect 22235 44693 22247 44696
rect 22189 44687 22247 44693
rect 22830 44684 22836 44696
rect 22888 44684 22894 44736
rect 23014 44724 23020 44736
rect 22975 44696 23020 44724
rect 23014 44684 23020 44696
rect 23072 44684 23078 44736
rect 23658 44724 23664 44736
rect 23619 44696 23664 44724
rect 23658 44684 23664 44696
rect 23716 44684 23722 44736
rect 26970 44684 26976 44736
rect 27028 44724 27034 44736
rect 27157 44727 27215 44733
rect 27157 44724 27169 44727
rect 27028 44696 27169 44724
rect 27028 44684 27034 44696
rect 27157 44693 27169 44696
rect 27203 44693 27215 44727
rect 27157 44687 27215 44693
rect 1104 44634 38824 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 38824 44634
rect 1104 44560 38824 44582
rect 20070 44480 20076 44532
rect 20128 44520 20134 44532
rect 20165 44523 20223 44529
rect 20165 44520 20177 44523
rect 20128 44492 20177 44520
rect 20128 44480 20134 44492
rect 20165 44489 20177 44492
rect 20211 44489 20223 44523
rect 21174 44520 21180 44532
rect 21135 44492 21180 44520
rect 20165 44483 20223 44489
rect 21174 44480 21180 44492
rect 21232 44480 21238 44532
rect 22189 44523 22247 44529
rect 22189 44489 22201 44523
rect 22235 44520 22247 44523
rect 23014 44520 23020 44532
rect 22235 44492 23020 44520
rect 22235 44489 22247 44492
rect 22189 44483 22247 44489
rect 23014 44480 23020 44492
rect 23072 44480 23078 44532
rect 27154 44520 27160 44532
rect 27115 44492 27160 44520
rect 27154 44480 27160 44492
rect 27212 44480 27218 44532
rect 36538 44480 36544 44532
rect 36596 44520 36602 44532
rect 37461 44523 37519 44529
rect 37461 44520 37473 44523
rect 36596 44492 37473 44520
rect 36596 44480 36602 44492
rect 37461 44489 37473 44492
rect 37507 44489 37519 44523
rect 37461 44483 37519 44489
rect 20714 44412 20720 44464
rect 20772 44452 20778 44464
rect 23324 44455 23382 44461
rect 20772 44424 21036 44452
rect 20772 44412 20778 44424
rect 18138 44384 18144 44396
rect 18099 44356 18144 44384
rect 18138 44344 18144 44356
rect 18196 44344 18202 44396
rect 18408 44387 18466 44393
rect 18408 44353 18420 44387
rect 18454 44384 18466 44387
rect 19242 44384 19248 44396
rect 18454 44356 19248 44384
rect 18454 44353 18466 44356
rect 18408 44347 18466 44353
rect 19242 44344 19248 44356
rect 19300 44344 19306 44396
rect 19978 44384 19984 44396
rect 19939 44356 19984 44384
rect 19978 44344 19984 44356
rect 20036 44344 20042 44396
rect 20898 44384 20904 44396
rect 20859 44356 20904 44384
rect 20898 44344 20904 44356
rect 20956 44344 20962 44396
rect 21008 44393 21036 44424
rect 23324 44421 23336 44455
rect 23370 44452 23382 44455
rect 23658 44452 23664 44464
rect 23370 44424 23664 44452
rect 23370 44421 23382 44424
rect 23324 44415 23382 44421
rect 23658 44412 23664 44424
rect 23716 44412 23722 44464
rect 20993 44387 21051 44393
rect 20993 44353 21005 44387
rect 21039 44384 21051 44387
rect 21450 44384 21456 44396
rect 21039 44356 21456 44384
rect 21039 44353 21051 44356
rect 20993 44347 21051 44353
rect 21450 44344 21456 44356
rect 21508 44344 21514 44396
rect 23566 44384 23572 44396
rect 23479 44356 23572 44384
rect 23566 44344 23572 44356
rect 23624 44384 23630 44396
rect 23934 44384 23940 44396
rect 23624 44356 23940 44384
rect 23624 44344 23630 44356
rect 23934 44344 23940 44356
rect 23992 44384 23998 44396
rect 24762 44384 24768 44396
rect 23992 44356 24768 44384
rect 23992 44344 23998 44356
rect 24762 44344 24768 44356
rect 24820 44344 24826 44396
rect 26050 44384 26056 44396
rect 26011 44356 26056 44384
rect 26050 44344 26056 44356
rect 26108 44344 26114 44396
rect 26970 44384 26976 44396
rect 26931 44356 26976 44384
rect 26970 44344 26976 44356
rect 27028 44344 27034 44396
rect 27798 44384 27804 44396
rect 27759 44356 27804 44384
rect 27798 44344 27804 44356
rect 27856 44344 27862 44396
rect 29914 44384 29920 44396
rect 29875 44356 29920 44384
rect 29914 44344 29920 44356
rect 29972 44344 29978 44396
rect 36722 44384 36728 44396
rect 36683 44356 36728 44384
rect 36722 44344 36728 44356
rect 36780 44344 36786 44396
rect 37366 44384 37372 44396
rect 37327 44356 37372 44384
rect 37366 44344 37372 44356
rect 37424 44344 37430 44396
rect 26234 44276 26240 44328
rect 26292 44316 26298 44328
rect 26292 44288 26337 44316
rect 26292 44276 26298 44288
rect 29270 44208 29276 44260
rect 29328 44248 29334 44260
rect 37366 44248 37372 44260
rect 29328 44220 37372 44248
rect 29328 44208 29334 44220
rect 37366 44208 37372 44220
rect 37424 44208 37430 44260
rect 19426 44140 19432 44192
rect 19484 44180 19490 44192
rect 19521 44183 19579 44189
rect 19521 44180 19533 44183
rect 19484 44152 19533 44180
rect 19484 44140 19490 44152
rect 19521 44149 19533 44152
rect 19567 44180 19579 44183
rect 20254 44180 20260 44192
rect 19567 44152 20260 44180
rect 19567 44149 19579 44152
rect 19521 44143 19579 44149
rect 20254 44140 20260 44152
rect 20312 44140 20318 44192
rect 25869 44183 25927 44189
rect 25869 44149 25881 44183
rect 25915 44180 25927 44183
rect 25958 44180 25964 44192
rect 25915 44152 25964 44180
rect 25915 44149 25927 44152
rect 25869 44143 25927 44149
rect 25958 44140 25964 44152
rect 26016 44140 26022 44192
rect 27982 44180 27988 44192
rect 27943 44152 27988 44180
rect 27982 44140 27988 44152
rect 28040 44140 28046 44192
rect 29733 44183 29791 44189
rect 29733 44149 29745 44183
rect 29779 44180 29791 44183
rect 29822 44180 29828 44192
rect 29779 44152 29828 44180
rect 29779 44149 29791 44152
rect 29733 44143 29791 44149
rect 29822 44140 29828 44152
rect 29880 44140 29886 44192
rect 1104 44090 38824 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 38824 44090
rect 1104 44016 38824 44038
rect 19242 43976 19248 43988
rect 19203 43948 19248 43976
rect 19242 43936 19248 43948
rect 19300 43936 19306 43988
rect 22005 43979 22063 43985
rect 22005 43945 22017 43979
rect 22051 43976 22063 43979
rect 23106 43976 23112 43988
rect 22051 43948 23112 43976
rect 22051 43945 22063 43948
rect 22005 43939 22063 43945
rect 23106 43936 23112 43948
rect 23164 43936 23170 43988
rect 25774 43976 25780 43988
rect 25735 43948 25780 43976
rect 25774 43936 25780 43948
rect 25832 43936 25838 43988
rect 27157 43979 27215 43985
rect 27157 43945 27169 43979
rect 27203 43976 27215 43979
rect 27798 43976 27804 43988
rect 27203 43948 27804 43976
rect 27203 43945 27215 43948
rect 27157 43939 27215 43945
rect 27798 43936 27804 43948
rect 27856 43936 27862 43988
rect 21637 43843 21695 43849
rect 6886 43812 16620 43840
rect 5442 43732 5448 43784
rect 5500 43772 5506 43784
rect 6886 43772 6914 43812
rect 16592 43781 16620 43812
rect 21637 43809 21649 43843
rect 21683 43840 21695 43843
rect 22094 43840 22100 43852
rect 21683 43812 22100 43840
rect 21683 43809 21695 43812
rect 21637 43803 21695 43809
rect 22094 43800 22100 43812
rect 22152 43800 22158 43852
rect 26050 43800 26056 43852
rect 26108 43840 26114 43852
rect 38102 43840 38108 43852
rect 26108 43812 27016 43840
rect 38063 43812 38108 43840
rect 26108 43800 26114 43812
rect 5500 43744 6914 43772
rect 16485 43775 16543 43781
rect 5500 43732 5506 43744
rect 16485 43741 16497 43775
rect 16531 43741 16543 43775
rect 16485 43735 16543 43741
rect 16577 43775 16635 43781
rect 16577 43741 16589 43775
rect 16623 43741 16635 43775
rect 16577 43735 16635 43741
rect 16761 43775 16819 43781
rect 16761 43741 16773 43775
rect 16807 43772 16819 43775
rect 17405 43775 17463 43781
rect 17405 43772 17417 43775
rect 16807 43744 17417 43772
rect 16807 43741 16819 43744
rect 16761 43735 16819 43741
rect 17405 43741 17417 43744
rect 17451 43741 17463 43775
rect 19426 43772 19432 43784
rect 19387 43744 19432 43772
rect 17405 43735 17463 43741
rect 16500 43704 16528 43735
rect 19426 43732 19432 43744
rect 19484 43732 19490 43784
rect 21450 43732 21456 43784
rect 21508 43772 21514 43784
rect 21821 43775 21879 43781
rect 21821 43772 21833 43775
rect 21508 43744 21833 43772
rect 21508 43732 21514 43744
rect 21821 43741 21833 43744
rect 21867 43741 21879 43775
rect 21821 43735 21879 43741
rect 25317 43775 25375 43781
rect 25317 43741 25329 43775
rect 25363 43772 25375 43775
rect 25774 43772 25780 43784
rect 25363 43744 25780 43772
rect 25363 43741 25375 43744
rect 25317 43735 25375 43741
rect 25774 43732 25780 43744
rect 25832 43732 25838 43784
rect 25958 43772 25964 43784
rect 25919 43744 25964 43772
rect 25958 43732 25964 43744
rect 26016 43732 26022 43784
rect 26878 43772 26884 43784
rect 26839 43744 26884 43772
rect 26878 43732 26884 43744
rect 26936 43732 26942 43784
rect 26988 43781 27016 43812
rect 38102 43800 38108 43812
rect 38160 43800 38166 43852
rect 26973 43775 27031 43781
rect 26973 43741 26985 43775
rect 27019 43741 27031 43775
rect 27614 43772 27620 43784
rect 27575 43744 27620 43772
rect 26973 43735 27031 43741
rect 27614 43732 27620 43744
rect 27672 43772 27678 43784
rect 28350 43772 28356 43784
rect 27672 43744 28356 43772
rect 27672 43732 27678 43744
rect 28350 43732 28356 43744
rect 28408 43772 28414 43784
rect 29822 43781 29828 43784
rect 29549 43775 29607 43781
rect 29549 43772 29561 43775
rect 28408 43744 29561 43772
rect 28408 43732 28414 43744
rect 29549 43741 29561 43744
rect 29595 43741 29607 43775
rect 29816 43772 29828 43781
rect 29783 43744 29828 43772
rect 29549 43735 29607 43741
rect 29816 43735 29828 43744
rect 29822 43732 29828 43735
rect 29880 43732 29886 43784
rect 36262 43772 36268 43784
rect 36223 43744 36268 43772
rect 36262 43732 36268 43744
rect 36320 43732 36326 43784
rect 16666 43704 16672 43716
rect 16500 43676 16672 43704
rect 16666 43664 16672 43676
rect 16724 43664 16730 43716
rect 27884 43707 27942 43713
rect 27884 43673 27896 43707
rect 27930 43704 27942 43707
rect 27982 43704 27988 43716
rect 27930 43676 27988 43704
rect 27930 43673 27942 43676
rect 27884 43667 27942 43673
rect 27982 43664 27988 43676
rect 28040 43664 28046 43716
rect 36449 43707 36507 43713
rect 36449 43673 36461 43707
rect 36495 43704 36507 43707
rect 37458 43704 37464 43716
rect 36495 43676 37464 43704
rect 36495 43673 36507 43676
rect 36449 43667 36507 43673
rect 37458 43664 37464 43676
rect 37516 43664 37522 43716
rect 17218 43636 17224 43648
rect 17179 43608 17224 43636
rect 17218 43596 17224 43608
rect 17276 43596 17282 43648
rect 25130 43636 25136 43648
rect 25091 43608 25136 43636
rect 25130 43596 25136 43608
rect 25188 43596 25194 43648
rect 28997 43639 29055 43645
rect 28997 43605 29009 43639
rect 29043 43636 29055 43639
rect 29546 43636 29552 43648
rect 29043 43608 29552 43636
rect 29043 43605 29055 43608
rect 28997 43599 29055 43605
rect 29546 43596 29552 43608
rect 29604 43596 29610 43648
rect 30926 43636 30932 43648
rect 30887 43608 30932 43636
rect 30926 43596 30932 43608
rect 30984 43596 30990 43648
rect 1104 43546 38824 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 38824 43546
rect 1104 43472 38824 43494
rect 19426 43432 19432 43444
rect 19387 43404 19432 43432
rect 19426 43392 19432 43404
rect 19484 43392 19490 43444
rect 25774 43432 25780 43444
rect 25735 43404 25780 43432
rect 25774 43392 25780 43404
rect 25832 43392 25838 43444
rect 26878 43392 26884 43444
rect 26936 43432 26942 43444
rect 27249 43435 27307 43441
rect 27249 43432 27261 43435
rect 26936 43404 27261 43432
rect 26936 43392 26942 43404
rect 27249 43401 27261 43404
rect 27295 43401 27307 43435
rect 27249 43395 27307 43401
rect 27338 43392 27344 43444
rect 27396 43432 27402 43444
rect 29914 43432 29920 43444
rect 27396 43404 27441 43432
rect 29875 43404 29920 43432
rect 27396 43392 27402 43404
rect 29914 43392 29920 43404
rect 29972 43392 29978 43444
rect 37458 43432 37464 43444
rect 37419 43404 37464 43432
rect 37458 43392 37464 43404
rect 37516 43392 37522 43444
rect 17028 43367 17086 43373
rect 17028 43333 17040 43367
rect 17074 43364 17086 43367
rect 17218 43364 17224 43376
rect 17074 43336 17224 43364
rect 17074 43333 17086 43336
rect 17028 43327 17086 43333
rect 17218 43324 17224 43336
rect 17276 43324 17282 43376
rect 19889 43367 19947 43373
rect 19889 43364 19901 43367
rect 19168 43336 19901 43364
rect 19168 43305 19196 43336
rect 19889 43333 19901 43336
rect 19935 43364 19947 43367
rect 19978 43364 19984 43376
rect 19935 43336 19984 43364
rect 19935 43333 19947 43336
rect 19889 43327 19947 43333
rect 19978 43324 19984 43336
rect 20036 43324 20042 43376
rect 26050 43364 26056 43376
rect 22940 43336 26056 43364
rect 19153 43299 19211 43305
rect 19153 43265 19165 43299
rect 19199 43265 19211 43299
rect 19153 43259 19211 43265
rect 19245 43299 19303 43305
rect 19245 43265 19257 43299
rect 19291 43265 19303 43299
rect 20162 43296 20168 43308
rect 20123 43268 20168 43296
rect 19245 43259 19303 43265
rect 16574 43188 16580 43240
rect 16632 43228 16638 43240
rect 16761 43231 16819 43237
rect 16761 43228 16773 43231
rect 16632 43200 16773 43228
rect 16632 43188 16638 43200
rect 16761 43197 16773 43200
rect 16807 43197 16819 43231
rect 16761 43191 16819 43197
rect 19260 43160 19288 43259
rect 20162 43256 20168 43268
rect 20220 43256 20226 43308
rect 22940 43305 22968 43336
rect 22925 43299 22983 43305
rect 22925 43265 22937 43299
rect 22971 43265 22983 43299
rect 23934 43296 23940 43308
rect 23895 43268 23940 43296
rect 22925 43259 22983 43265
rect 23934 43256 23940 43268
rect 23992 43256 23998 43308
rect 24026 43256 24032 43308
rect 24084 43296 24090 43308
rect 25976 43305 26004 43336
rect 26050 43324 26056 43336
rect 26108 43324 26114 43376
rect 24193 43299 24251 43305
rect 24193 43296 24205 43299
rect 24084 43268 24205 43296
rect 24084 43256 24090 43268
rect 24193 43265 24205 43268
rect 24239 43265 24251 43299
rect 24193 43259 24251 43265
rect 25961 43299 26019 43305
rect 25961 43265 25973 43299
rect 26007 43265 26019 43299
rect 25961 43259 26019 43265
rect 27062 43256 27068 43308
rect 27120 43296 27126 43308
rect 27157 43299 27215 43305
rect 27157 43296 27169 43299
rect 27120 43268 27169 43296
rect 27120 43256 27126 43268
rect 27157 43265 27169 43268
rect 27203 43265 27215 43299
rect 29546 43296 29552 43308
rect 29507 43268 29552 43296
rect 27157 43259 27215 43265
rect 29546 43256 29552 43268
rect 29604 43256 29610 43308
rect 29733 43299 29791 43305
rect 29733 43265 29745 43299
rect 29779 43296 29791 43299
rect 30282 43296 30288 43308
rect 29779 43268 30288 43296
rect 29779 43265 29791 43268
rect 29733 43259 29791 43265
rect 30282 43256 30288 43268
rect 30340 43256 30346 43308
rect 31110 43296 31116 43308
rect 31071 43268 31116 43296
rect 31110 43256 31116 43268
rect 31168 43256 31174 43308
rect 35802 43256 35808 43308
rect 35860 43296 35866 43308
rect 36081 43299 36139 43305
rect 36081 43296 36093 43299
rect 35860 43268 36093 43296
rect 35860 43256 35866 43268
rect 36081 43265 36093 43268
rect 36127 43265 36139 43299
rect 36081 43259 36139 43265
rect 36262 43256 36268 43308
rect 36320 43296 36326 43308
rect 36541 43299 36599 43305
rect 36541 43296 36553 43299
rect 36320 43268 36553 43296
rect 36320 43256 36326 43268
rect 36541 43265 36553 43268
rect 36587 43265 36599 43299
rect 36541 43259 36599 43265
rect 37369 43299 37427 43305
rect 37369 43265 37381 43299
rect 37415 43296 37427 43299
rect 37826 43296 37832 43308
rect 37415 43268 37832 43296
rect 37415 43265 37427 43268
rect 37369 43259 37427 43265
rect 37826 43256 37832 43268
rect 37884 43256 37890 43308
rect 20073 43231 20131 43237
rect 20073 43197 20085 43231
rect 20119 43228 20131 43231
rect 20254 43228 20260 43240
rect 20119 43200 20260 43228
rect 20119 43197 20131 43200
rect 20073 43191 20131 43197
rect 20254 43188 20260 43200
rect 20312 43188 20318 43240
rect 21174 43188 21180 43240
rect 21232 43228 21238 43240
rect 22649 43231 22707 43237
rect 22649 43228 22661 43231
rect 21232 43200 22661 43228
rect 21232 43188 21238 43200
rect 22649 43197 22661 43200
rect 22695 43197 22707 43231
rect 26145 43231 26203 43237
rect 26145 43228 26157 43231
rect 22649 43191 22707 43197
rect 25332 43200 26157 43228
rect 21450 43160 21456 43172
rect 19260 43132 21456 43160
rect 21450 43120 21456 43132
rect 21508 43120 21514 43172
rect 25332 43169 25360 43200
rect 26145 43197 26157 43200
rect 26191 43228 26203 43231
rect 27080 43228 27108 43256
rect 26191 43200 27108 43228
rect 26191 43197 26203 43200
rect 26145 43191 26203 43197
rect 25317 43163 25375 43169
rect 25317 43129 25329 43163
rect 25363 43129 25375 43163
rect 25317 43123 25375 43129
rect 26234 43120 26240 43172
rect 26292 43160 26298 43172
rect 26970 43160 26976 43172
rect 26292 43132 26976 43160
rect 26292 43120 26298 43132
rect 26970 43120 26976 43132
rect 27028 43120 27034 43172
rect 1578 43092 1584 43104
rect 1539 43064 1584 43092
rect 1578 43052 1584 43064
rect 1636 43052 1642 43104
rect 2038 43052 2044 43104
rect 2096 43092 2102 43104
rect 2225 43095 2283 43101
rect 2225 43092 2237 43095
rect 2096 43064 2237 43092
rect 2096 43052 2102 43064
rect 2225 43061 2237 43064
rect 2271 43061 2283 43095
rect 2225 43055 2283 43061
rect 18141 43095 18199 43101
rect 18141 43061 18153 43095
rect 18187 43092 18199 43095
rect 18230 43092 18236 43104
rect 18187 43064 18236 43092
rect 18187 43061 18199 43064
rect 18141 43055 18199 43061
rect 18230 43052 18236 43064
rect 18288 43092 18294 43104
rect 19242 43092 19248 43104
rect 18288 43064 19248 43092
rect 18288 43052 18294 43064
rect 19242 43052 19248 43064
rect 19300 43092 19306 43104
rect 19889 43095 19947 43101
rect 19889 43092 19901 43095
rect 19300 43064 19901 43092
rect 19300 43052 19306 43064
rect 19889 43061 19901 43064
rect 19935 43061 19947 43095
rect 19889 43055 19947 43061
rect 20349 43095 20407 43101
rect 20349 43061 20361 43095
rect 20395 43092 20407 43095
rect 21266 43092 21272 43104
rect 20395 43064 21272 43092
rect 20395 43061 20407 43064
rect 20349 43055 20407 43061
rect 21266 43052 21272 43064
rect 21324 43052 21330 43104
rect 27154 43052 27160 43104
rect 27212 43092 27218 43104
rect 27525 43095 27583 43101
rect 27525 43092 27537 43095
rect 27212 43064 27537 43092
rect 27212 43052 27218 43064
rect 27525 43061 27537 43064
rect 27571 43061 27583 43095
rect 27525 43055 27583 43061
rect 31297 43095 31355 43101
rect 31297 43061 31309 43095
rect 31343 43092 31355 43095
rect 31938 43092 31944 43104
rect 31343 43064 31944 43092
rect 31343 43061 31355 43064
rect 31297 43055 31355 43061
rect 31938 43052 31944 43064
rect 31996 43052 32002 43104
rect 35894 43052 35900 43104
rect 35952 43092 35958 43104
rect 35952 43064 35997 43092
rect 35952 43052 35958 43064
rect 1104 43002 38824 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 38824 43002
rect 1104 42928 38824 42950
rect 22646 42848 22652 42900
rect 22704 42888 22710 42900
rect 22704 42860 25820 42888
rect 22704 42848 22710 42860
rect 19981 42823 20039 42829
rect 19981 42789 19993 42823
rect 20027 42820 20039 42823
rect 20162 42820 20168 42832
rect 20027 42792 20168 42820
rect 20027 42789 20039 42792
rect 19981 42783 20039 42789
rect 20162 42780 20168 42792
rect 20220 42780 20226 42832
rect 25792 42820 25820 42860
rect 26234 42848 26240 42900
rect 26292 42888 26298 42900
rect 27062 42888 27068 42900
rect 26292 42860 26337 42888
rect 27023 42860 27068 42888
rect 26292 42848 26298 42860
rect 27062 42848 27068 42860
rect 27120 42848 27126 42900
rect 37826 42888 37832 42900
rect 31036 42860 37832 42888
rect 31036 42820 31064 42860
rect 37826 42848 37832 42860
rect 37884 42848 37890 42900
rect 25792 42792 31064 42820
rect 1397 42755 1455 42761
rect 1397 42721 1409 42755
rect 1443 42752 1455 42755
rect 1578 42752 1584 42764
rect 1443 42724 1584 42752
rect 1443 42721 1455 42724
rect 1397 42715 1455 42721
rect 1578 42712 1584 42724
rect 1636 42712 1642 42764
rect 2774 42752 2780 42764
rect 2735 42724 2780 42752
rect 2774 42712 2780 42724
rect 2832 42712 2838 42764
rect 16666 42712 16672 42764
rect 16724 42752 16730 42764
rect 17221 42755 17279 42761
rect 17221 42752 17233 42755
rect 16724 42724 17233 42752
rect 16724 42712 16730 42724
rect 17221 42721 17233 42724
rect 17267 42752 17279 42755
rect 23474 42752 23480 42764
rect 17267 42724 23480 42752
rect 17267 42721 17279 42724
rect 17221 42715 17279 42721
rect 23474 42712 23480 42724
rect 23532 42712 23538 42764
rect 23566 42712 23572 42764
rect 23624 42752 23630 42764
rect 23934 42752 23940 42764
rect 23624 42724 23940 42752
rect 23624 42712 23630 42724
rect 23934 42712 23940 42724
rect 23992 42752 23998 42764
rect 24857 42755 24915 42761
rect 24857 42752 24869 42755
rect 23992 42724 24869 42752
rect 23992 42712 23998 42724
rect 24857 42721 24869 42724
rect 24903 42721 24915 42755
rect 26878 42752 26884 42764
rect 26839 42724 26884 42752
rect 24857 42715 24915 42721
rect 26878 42712 26884 42724
rect 26936 42712 26942 42764
rect 30101 42755 30159 42761
rect 30101 42721 30113 42755
rect 30147 42752 30159 42755
rect 30374 42752 30380 42764
rect 30147 42724 30380 42752
rect 30147 42721 30159 42724
rect 30101 42715 30159 42721
rect 30374 42712 30380 42724
rect 30432 42752 30438 42764
rect 30926 42752 30932 42764
rect 30432 42724 30932 42752
rect 30432 42712 30438 42724
rect 30926 42712 30932 42724
rect 30984 42712 30990 42764
rect 16209 42687 16267 42693
rect 16209 42653 16221 42687
rect 16255 42684 16267 42687
rect 16853 42687 16911 42693
rect 16853 42684 16865 42687
rect 16255 42656 16865 42684
rect 16255 42653 16267 42656
rect 16209 42647 16267 42653
rect 16853 42653 16865 42656
rect 16899 42653 16911 42687
rect 16853 42647 16911 42653
rect 17037 42687 17095 42693
rect 17037 42653 17049 42687
rect 17083 42653 17095 42687
rect 17037 42647 17095 42653
rect 1578 42616 1584 42628
rect 1539 42588 1584 42616
rect 1578 42576 1584 42588
rect 1636 42576 1642 42628
rect 17052 42616 17080 42647
rect 18598 42644 18604 42696
rect 18656 42684 18662 42696
rect 18693 42687 18751 42693
rect 18693 42684 18705 42687
rect 18656 42656 18705 42684
rect 18656 42644 18662 42656
rect 18693 42653 18705 42656
rect 18739 42653 18751 42687
rect 20806 42684 20812 42696
rect 18693 42647 18751 42653
rect 18800 42656 20812 42684
rect 18800 42616 18828 42656
rect 20806 42644 20812 42656
rect 20864 42644 20870 42696
rect 21174 42684 21180 42696
rect 21135 42656 21180 42684
rect 21174 42644 21180 42656
rect 21232 42644 21238 42696
rect 21450 42684 21456 42696
rect 21411 42656 21456 42684
rect 21450 42644 21456 42656
rect 21508 42644 21514 42696
rect 22186 42644 22192 42696
rect 22244 42684 22250 42696
rect 25130 42693 25136 42696
rect 22465 42687 22523 42693
rect 22465 42684 22477 42687
rect 22244 42656 22477 42684
rect 22244 42644 22250 42656
rect 22465 42653 22477 42656
rect 22511 42653 22523 42687
rect 22465 42647 22523 42653
rect 23661 42687 23719 42693
rect 23661 42653 23673 42687
rect 23707 42653 23719 42687
rect 25124 42684 25136 42693
rect 25091 42656 25136 42684
rect 23661 42647 23719 42653
rect 25124 42647 25136 42656
rect 17052 42588 18828 42616
rect 19978 42576 19984 42628
rect 20036 42616 20042 42628
rect 20349 42619 20407 42625
rect 20349 42616 20361 42619
rect 20036 42588 20361 42616
rect 20036 42576 20042 42588
rect 20349 42585 20361 42588
rect 20395 42585 20407 42619
rect 20349 42579 20407 42585
rect 21266 42576 21272 42628
rect 21324 42616 21330 42628
rect 22649 42619 22707 42625
rect 22649 42616 22661 42619
rect 21324 42588 22661 42616
rect 21324 42576 21330 42588
rect 22649 42585 22661 42588
rect 22695 42585 22707 42619
rect 23676 42616 23704 42647
rect 25130 42644 25136 42647
rect 25188 42644 25194 42696
rect 26970 42644 26976 42696
rect 27028 42684 27034 42696
rect 27065 42687 27123 42693
rect 27065 42684 27077 42687
rect 27028 42656 27077 42684
rect 27028 42644 27034 42656
rect 27065 42653 27077 42656
rect 27111 42653 27123 42687
rect 27338 42684 27344 42696
rect 27065 42647 27123 42653
rect 27172 42656 27344 42684
rect 23934 42616 23940 42628
rect 23676 42588 23940 42616
rect 22649 42579 22707 42585
rect 23934 42576 23940 42588
rect 23992 42576 23998 42628
rect 26789 42619 26847 42625
rect 26789 42585 26801 42619
rect 26835 42616 26847 42619
rect 27172 42616 27200 42656
rect 27338 42644 27344 42656
rect 27396 42644 27402 42696
rect 29733 42687 29791 42693
rect 29733 42653 29745 42687
rect 29779 42684 29791 42687
rect 29914 42684 29920 42696
rect 29779 42656 29920 42684
rect 29779 42653 29791 42656
rect 29733 42647 29791 42653
rect 29914 42644 29920 42656
rect 29972 42684 29978 42696
rect 29972 42656 30880 42684
rect 29972 42644 29978 42656
rect 27893 42619 27951 42625
rect 27893 42616 27905 42619
rect 26835 42588 27200 42616
rect 27264 42588 27905 42616
rect 26835 42585 26847 42588
rect 26789 42579 26847 42585
rect 16393 42551 16451 42557
rect 16393 42517 16405 42551
rect 16439 42548 16451 42551
rect 16482 42548 16488 42560
rect 16439 42520 16488 42548
rect 16439 42517 16451 42520
rect 16393 42511 16451 42517
rect 16482 42508 16488 42520
rect 16540 42508 16546 42560
rect 18322 42508 18328 42560
rect 18380 42548 18386 42560
rect 18509 42551 18567 42557
rect 18509 42548 18521 42551
rect 18380 42520 18521 42548
rect 18380 42508 18386 42520
rect 18509 42517 18521 42520
rect 18555 42517 18567 42551
rect 18509 42511 18567 42517
rect 19242 42508 19248 42560
rect 19300 42548 19306 42560
rect 20165 42551 20223 42557
rect 20165 42548 20177 42551
rect 19300 42520 20177 42548
rect 19300 42508 19306 42520
rect 20165 42517 20177 42520
rect 20211 42517 20223 42551
rect 20165 42511 20223 42517
rect 20254 42508 20260 42560
rect 20312 42548 20318 42560
rect 20533 42551 20591 42557
rect 20312 42520 20357 42548
rect 20312 42508 20318 42520
rect 20533 42517 20545 42551
rect 20579 42548 20591 42551
rect 22278 42548 22284 42560
rect 20579 42520 22284 42548
rect 20579 42517 20591 42520
rect 20533 42511 20591 42517
rect 22278 42508 22284 42520
rect 22336 42508 22342 42560
rect 22830 42548 22836 42560
rect 22791 42520 22836 42548
rect 22830 42508 22836 42520
rect 22888 42508 22894 42560
rect 23750 42508 23756 42560
rect 23808 42548 23814 42560
rect 27264 42557 27292 42588
rect 27893 42585 27905 42588
rect 27939 42585 27951 42619
rect 27893 42579 27951 42585
rect 28077 42619 28135 42625
rect 28077 42585 28089 42619
rect 28123 42616 28135 42619
rect 29362 42616 29368 42628
rect 28123 42588 29368 42616
rect 28123 42585 28135 42588
rect 28077 42579 28135 42585
rect 29362 42576 29368 42588
rect 29420 42576 29426 42628
rect 29825 42619 29883 42625
rect 29825 42585 29837 42619
rect 29871 42616 29883 42619
rect 30006 42616 30012 42628
rect 29871 42588 30012 42616
rect 29871 42585 29883 42588
rect 29825 42579 29883 42585
rect 30006 42576 30012 42588
rect 30064 42576 30070 42628
rect 23845 42551 23903 42557
rect 23845 42548 23857 42551
rect 23808 42520 23857 42548
rect 23808 42508 23814 42520
rect 23845 42517 23857 42520
rect 23891 42517 23903 42551
rect 23845 42511 23903 42517
rect 27249 42551 27307 42557
rect 27249 42517 27261 42551
rect 27295 42517 27307 42551
rect 27706 42548 27712 42560
rect 27667 42520 27712 42548
rect 27249 42511 27307 42517
rect 27706 42508 27712 42520
rect 27764 42508 27770 42560
rect 27798 42508 27804 42560
rect 27856 42548 27862 42560
rect 29549 42551 29607 42557
rect 29549 42548 29561 42551
rect 27856 42520 29561 42548
rect 27856 42508 27862 42520
rect 29549 42517 29561 42520
rect 29595 42517 29607 42551
rect 29549 42511 29607 42517
rect 29638 42508 29644 42560
rect 29696 42548 29702 42560
rect 30852 42557 30880 42656
rect 31938 42644 31944 42696
rect 31996 42693 32002 42696
rect 31996 42684 32008 42693
rect 32217 42687 32275 42693
rect 31996 42656 32041 42684
rect 31996 42647 32008 42656
rect 32217 42653 32229 42687
rect 32263 42684 32275 42687
rect 33042 42684 33048 42696
rect 32263 42656 33048 42684
rect 32263 42653 32275 42656
rect 32217 42647 32275 42653
rect 31996 42644 32002 42647
rect 33042 42644 33048 42656
rect 33100 42644 33106 42696
rect 36262 42684 36268 42696
rect 36223 42656 36268 42684
rect 36262 42644 36268 42656
rect 36320 42644 36326 42696
rect 36446 42616 36452 42628
rect 36407 42588 36452 42616
rect 36446 42576 36452 42588
rect 36504 42576 36510 42628
rect 38102 42616 38108 42628
rect 38063 42588 38108 42616
rect 38102 42576 38108 42588
rect 38160 42576 38166 42628
rect 29917 42551 29975 42557
rect 29917 42548 29929 42551
rect 29696 42520 29929 42548
rect 29696 42508 29702 42520
rect 29917 42517 29929 42520
rect 29963 42517 29975 42551
rect 29917 42511 29975 42517
rect 30837 42551 30895 42557
rect 30837 42517 30849 42551
rect 30883 42517 30895 42551
rect 30837 42511 30895 42517
rect 1104 42458 38824 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 38824 42458
rect 1104 42384 38824 42406
rect 1489 42347 1547 42353
rect 1489 42313 1501 42347
rect 1535 42344 1547 42347
rect 1578 42344 1584 42356
rect 1535 42316 1584 42344
rect 1535 42313 1547 42316
rect 1489 42307 1547 42313
rect 1578 42304 1584 42316
rect 1636 42304 1642 42356
rect 19429 42347 19487 42353
rect 19429 42313 19441 42347
rect 19475 42344 19487 42347
rect 20162 42344 20168 42356
rect 19475 42316 20168 42344
rect 19475 42313 19487 42316
rect 19429 42307 19487 42313
rect 20162 42304 20168 42316
rect 20220 42304 20226 42356
rect 23290 42344 23296 42356
rect 22480 42316 23296 42344
rect 22480 42285 22508 42316
rect 23290 42304 23296 42316
rect 23348 42304 23354 42356
rect 23937 42347 23995 42353
rect 23937 42313 23949 42347
rect 23983 42344 23995 42347
rect 24026 42344 24032 42356
rect 23983 42316 24032 42344
rect 23983 42313 23995 42316
rect 23937 42307 23995 42313
rect 24026 42304 24032 42316
rect 24084 42304 24090 42356
rect 27798 42344 27804 42356
rect 27264 42316 27804 42344
rect 27264 42285 27292 42316
rect 27798 42304 27804 42316
rect 27856 42304 27862 42356
rect 29362 42344 29368 42356
rect 29323 42316 29368 42344
rect 29362 42304 29368 42316
rect 29420 42304 29426 42356
rect 30745 42347 30803 42353
rect 30745 42313 30757 42347
rect 30791 42344 30803 42347
rect 31110 42344 31116 42356
rect 30791 42316 31116 42344
rect 30791 42313 30803 42316
rect 30745 42307 30803 42313
rect 31110 42304 31116 42316
rect 31168 42304 31174 42356
rect 36446 42304 36452 42356
rect 36504 42344 36510 42356
rect 37553 42347 37611 42353
rect 37553 42344 37565 42347
rect 36504 42316 37565 42344
rect 36504 42304 36510 42316
rect 37553 42313 37565 42316
rect 37599 42313 37611 42347
rect 37553 42307 37611 42313
rect 22465 42279 22523 42285
rect 18064 42248 21312 42276
rect 1581 42211 1639 42217
rect 1581 42177 1593 42211
rect 1627 42177 1639 42211
rect 2038 42208 2044 42220
rect 1999 42180 2044 42208
rect 1581 42171 1639 42177
rect 1596 42072 1624 42171
rect 2038 42168 2044 42180
rect 2096 42168 2102 42220
rect 9674 42208 9680 42220
rect 9635 42180 9680 42208
rect 9674 42168 9680 42180
rect 9732 42168 9738 42220
rect 16574 42168 16580 42220
rect 16632 42208 16638 42220
rect 18064 42217 18092 42248
rect 18322 42217 18328 42220
rect 18049 42211 18107 42217
rect 18049 42208 18061 42211
rect 16632 42180 18061 42208
rect 16632 42168 16638 42180
rect 18049 42177 18061 42180
rect 18095 42177 18107 42211
rect 18316 42208 18328 42217
rect 18283 42180 18328 42208
rect 18049 42171 18107 42177
rect 18316 42171 18328 42180
rect 18322 42168 18328 42171
rect 18380 42168 18386 42220
rect 20990 42208 20996 42220
rect 21048 42217 21054 42220
rect 20960 42180 20996 42208
rect 20990 42168 20996 42180
rect 21048 42171 21060 42217
rect 21048 42168 21054 42171
rect 21284 42152 21312 42248
rect 22465 42245 22477 42279
rect 22511 42245 22523 42279
rect 22465 42239 22523 42245
rect 27249 42279 27307 42285
rect 27249 42245 27261 42279
rect 27295 42245 27307 42279
rect 27249 42239 27307 42245
rect 27479 42279 27537 42285
rect 27479 42245 27491 42279
rect 27525 42276 27537 42279
rect 27706 42276 27712 42288
rect 27525 42248 27712 42276
rect 27525 42245 27537 42248
rect 27479 42239 27537 42245
rect 27706 42236 27712 42248
rect 27764 42236 27770 42288
rect 29825 42279 29883 42285
rect 29825 42245 29837 42279
rect 29871 42276 29883 42279
rect 29914 42276 29920 42288
rect 29871 42248 29920 42276
rect 29871 42245 29883 42248
rect 29825 42239 29883 42245
rect 29914 42236 29920 42248
rect 29972 42236 29978 42288
rect 22278 42208 22284 42220
rect 22239 42180 22284 42208
rect 22278 42168 22284 42180
rect 22336 42168 22342 42220
rect 22370 42168 22376 42220
rect 22428 42208 22434 42220
rect 22603 42211 22661 42217
rect 22428 42180 22473 42208
rect 22428 42168 22434 42180
rect 22603 42177 22615 42211
rect 22649 42208 22661 42211
rect 22830 42208 22836 42220
rect 22649 42180 22836 42208
rect 22649 42177 22661 42180
rect 22603 42171 22661 42177
rect 22830 42168 22836 42180
rect 22888 42168 22894 42220
rect 23750 42208 23756 42220
rect 23711 42180 23756 42208
rect 23750 42168 23756 42180
rect 23808 42168 23814 42220
rect 27154 42208 27160 42220
rect 27115 42180 27160 42208
rect 27154 42168 27160 42180
rect 27212 42168 27218 42220
rect 27341 42211 27399 42217
rect 27341 42177 27353 42211
rect 27387 42177 27399 42211
rect 27341 42171 27399 42177
rect 29549 42211 29607 42217
rect 29549 42177 29561 42211
rect 29595 42208 29607 42211
rect 30374 42208 30380 42220
rect 29595 42180 30380 42208
rect 29595 42177 29607 42180
rect 29549 42171 29607 42177
rect 2225 42143 2283 42149
rect 2225 42109 2237 42143
rect 2271 42140 2283 42143
rect 2866 42140 2872 42152
rect 2271 42112 2872 42140
rect 2271 42109 2283 42112
rect 2225 42103 2283 42109
rect 2866 42100 2872 42112
rect 2924 42100 2930 42152
rect 2958 42100 2964 42152
rect 3016 42140 3022 42152
rect 10410 42140 10416 42152
rect 3016 42112 3061 42140
rect 10371 42112 10416 42140
rect 3016 42100 3022 42112
rect 10410 42100 10416 42112
rect 10468 42100 10474 42152
rect 21266 42140 21272 42152
rect 21227 42112 21272 42140
rect 21266 42100 21272 42112
rect 21324 42100 21330 42152
rect 22738 42140 22744 42152
rect 22699 42112 22744 42140
rect 22738 42100 22744 42112
rect 22796 42100 22802 42152
rect 23290 42100 23296 42152
rect 23348 42140 23354 42152
rect 27356 42140 27384 42171
rect 30374 42168 30380 42180
rect 30432 42168 30438 42220
rect 30466 42168 30472 42220
rect 30524 42208 30530 42220
rect 33870 42217 33876 42220
rect 30561 42211 30619 42217
rect 30561 42208 30573 42211
rect 30524 42180 30573 42208
rect 30524 42168 30530 42180
rect 30561 42177 30573 42180
rect 30607 42177 30619 42211
rect 30561 42171 30619 42177
rect 33864 42171 33876 42217
rect 33928 42208 33934 42220
rect 33928 42180 33964 42208
rect 33870 42168 33876 42171
rect 33928 42168 33934 42180
rect 36262 42168 36268 42220
rect 36320 42208 36326 42220
rect 36541 42211 36599 42217
rect 36541 42208 36553 42211
rect 36320 42180 36553 42208
rect 36320 42168 36326 42180
rect 36541 42177 36553 42180
rect 36587 42177 36599 42211
rect 36541 42171 36599 42177
rect 37366 42168 37372 42220
rect 37424 42208 37430 42220
rect 37461 42211 37519 42217
rect 37461 42208 37473 42211
rect 37424 42180 37473 42208
rect 37424 42168 37430 42180
rect 37461 42177 37473 42180
rect 37507 42177 37519 42211
rect 37461 42171 37519 42177
rect 23348 42112 27384 42140
rect 27617 42143 27675 42149
rect 23348 42100 23354 42112
rect 27617 42109 27629 42143
rect 27663 42140 27675 42143
rect 27706 42140 27712 42152
rect 27663 42112 27712 42140
rect 27663 42109 27675 42112
rect 27617 42103 27675 42109
rect 27706 42100 27712 42112
rect 27764 42100 27770 42152
rect 29733 42143 29791 42149
rect 29733 42109 29745 42143
rect 29779 42140 29791 42143
rect 30006 42140 30012 42152
rect 29779 42112 30012 42140
rect 29779 42109 29791 42112
rect 29733 42103 29791 42109
rect 30006 42100 30012 42112
rect 30064 42100 30070 42152
rect 33042 42100 33048 42152
rect 33100 42140 33106 42152
rect 33597 42143 33655 42149
rect 33597 42140 33609 42143
rect 33100 42112 33609 42140
rect 33100 42100 33106 42112
rect 33597 42109 33609 42112
rect 33643 42109 33655 42143
rect 33597 42103 33655 42109
rect 14458 42072 14464 42084
rect 1596 42044 14464 42072
rect 14458 42032 14464 42044
rect 14516 42032 14522 42084
rect 23842 42072 23848 42084
rect 18984 42044 20024 42072
rect 10410 41964 10416 42016
rect 10468 42004 10474 42016
rect 18984 42004 19012 42044
rect 19886 42004 19892 42016
rect 10468 41976 19012 42004
rect 19847 41976 19892 42004
rect 10468 41964 10474 41976
rect 19886 41964 19892 41976
rect 19944 41964 19950 42016
rect 19996 42004 20024 42044
rect 21284 42044 23848 42072
rect 21284 42004 21312 42044
rect 23842 42032 23848 42044
rect 23900 42032 23906 42084
rect 22094 42004 22100 42016
rect 19996 41976 21312 42004
rect 22055 41976 22100 42004
rect 22094 41964 22100 41976
rect 22152 41964 22158 42016
rect 26970 42004 26976 42016
rect 26931 41976 26976 42004
rect 26970 41964 26976 41976
rect 27028 41964 27034 42016
rect 29638 42004 29644 42016
rect 29599 41976 29644 42004
rect 29638 41964 29644 41976
rect 29696 41964 29702 42016
rect 34790 41964 34796 42016
rect 34848 42004 34854 42016
rect 34977 42007 35035 42013
rect 34977 42004 34989 42007
rect 34848 41976 34989 42004
rect 34848 41964 34854 41976
rect 34977 41973 34989 41976
rect 35023 41973 35035 42007
rect 34977 41967 35035 41973
rect 1104 41914 38824 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 38824 41914
rect 1104 41840 38824 41862
rect 2866 41800 2872 41812
rect 2827 41772 2872 41800
rect 2866 41760 2872 41772
rect 2924 41760 2930 41812
rect 18598 41800 18604 41812
rect 18559 41772 18604 41800
rect 18598 41760 18604 41772
rect 18656 41760 18662 41812
rect 20901 41803 20959 41809
rect 20901 41769 20913 41803
rect 20947 41800 20959 41803
rect 20990 41800 20996 41812
rect 20947 41772 20996 41800
rect 20947 41769 20959 41772
rect 20901 41763 20959 41769
rect 20990 41760 20996 41772
rect 21048 41760 21054 41812
rect 22738 41800 22744 41812
rect 22699 41772 22744 41800
rect 22738 41760 22744 41772
rect 22796 41760 22802 41812
rect 33870 41760 33876 41812
rect 33928 41800 33934 41812
rect 33965 41803 34023 41809
rect 33965 41800 33977 41803
rect 33928 41772 33977 41800
rect 33928 41760 33934 41772
rect 33965 41769 33977 41772
rect 34011 41769 34023 41803
rect 33965 41763 34023 41769
rect 10042 41664 10048 41676
rect 10003 41636 10048 41664
rect 10042 41624 10048 41636
rect 10100 41624 10106 41676
rect 18230 41664 18236 41676
rect 18191 41636 18236 41664
rect 18230 41624 18236 41636
rect 18288 41624 18294 41676
rect 19889 41667 19947 41673
rect 19889 41633 19901 41667
rect 19935 41664 19947 41667
rect 20162 41664 20168 41676
rect 19935 41636 20168 41664
rect 19935 41633 19947 41636
rect 19889 41627 19947 41633
rect 20162 41624 20168 41636
rect 20220 41624 20226 41676
rect 23474 41624 23480 41676
rect 23532 41664 23538 41676
rect 23842 41664 23848 41676
rect 23532 41636 23848 41664
rect 23532 41624 23538 41636
rect 23842 41624 23848 41636
rect 23900 41624 23906 41676
rect 29914 41664 29920 41676
rect 29875 41636 29920 41664
rect 29914 41624 29920 41636
rect 29972 41624 29978 41676
rect 31202 41664 31208 41676
rect 30852 41636 31208 41664
rect 1394 41596 1400 41608
rect 1355 41568 1400 41596
rect 1394 41556 1400 41568
rect 1452 41556 1458 41608
rect 2961 41599 3019 41605
rect 2961 41565 2973 41599
rect 3007 41596 3019 41599
rect 8846 41596 8852 41608
rect 3007 41568 8852 41596
rect 3007 41565 3019 41568
rect 2961 41559 3019 41565
rect 8846 41556 8852 41568
rect 8904 41556 8910 41608
rect 9674 41596 9680 41608
rect 9635 41568 9680 41596
rect 9674 41556 9680 41568
rect 9732 41556 9738 41608
rect 16482 41605 16488 41608
rect 16209 41599 16267 41605
rect 16209 41565 16221 41599
rect 16255 41565 16267 41599
rect 16209 41559 16267 41565
rect 16476 41559 16488 41605
rect 16540 41596 16546 41608
rect 18417 41599 18475 41605
rect 16540 41568 16576 41596
rect 16224 41528 16252 41559
rect 16482 41556 16488 41559
rect 16540 41556 16546 41568
rect 18417 41565 18429 41599
rect 18463 41596 18475 41599
rect 19426 41596 19432 41608
rect 18463 41568 19432 41596
rect 18463 41565 18475 41568
rect 18417 41559 18475 41565
rect 19426 41556 19432 41568
rect 19484 41556 19490 41608
rect 20073 41599 20131 41605
rect 20073 41565 20085 41599
rect 20119 41565 20131 41599
rect 20073 41559 20131 41565
rect 20257 41599 20315 41605
rect 20257 41565 20269 41599
rect 20303 41596 20315 41599
rect 20717 41599 20775 41605
rect 20717 41596 20729 41599
rect 20303 41568 20729 41596
rect 20303 41565 20315 41568
rect 20257 41559 20315 41565
rect 20717 41565 20729 41568
rect 20763 41565 20775 41599
rect 20717 41559 20775 41565
rect 22925 41599 22983 41605
rect 22925 41565 22937 41599
rect 22971 41596 22983 41599
rect 23658 41596 23664 41608
rect 22971 41568 23664 41596
rect 22971 41565 22983 41568
rect 22925 41559 22983 41565
rect 16574 41528 16580 41540
rect 16224 41500 16580 41528
rect 16574 41488 16580 41500
rect 16632 41488 16638 41540
rect 18046 41528 18052 41540
rect 17420 41500 18052 41528
rect 1581 41463 1639 41469
rect 1581 41429 1593 41463
rect 1627 41460 1639 41463
rect 8386 41460 8392 41472
rect 1627 41432 8392 41460
rect 1627 41429 1639 41432
rect 1581 41423 1639 41429
rect 8386 41420 8392 41432
rect 8444 41420 8450 41472
rect 10042 41420 10048 41472
rect 10100 41460 10106 41472
rect 17420 41460 17448 41500
rect 18046 41488 18052 41500
rect 18104 41528 18110 41540
rect 19242 41528 19248 41540
rect 18104 41500 19248 41528
rect 18104 41488 18110 41500
rect 19242 41488 19248 41500
rect 19300 41488 19306 41540
rect 20088 41528 20116 41559
rect 23658 41556 23664 41568
rect 23716 41556 23722 41608
rect 26970 41556 26976 41608
rect 27028 41596 27034 41608
rect 27442 41599 27500 41605
rect 27442 41596 27454 41599
rect 27028 41568 27454 41596
rect 27028 41556 27034 41568
rect 27442 41565 27454 41568
rect 27488 41565 27500 41599
rect 27442 41559 27500 41565
rect 27614 41556 27620 41608
rect 27672 41596 27678 41608
rect 27709 41599 27767 41605
rect 27709 41596 27721 41599
rect 27672 41568 27721 41596
rect 27672 41556 27678 41568
rect 27709 41565 27721 41568
rect 27755 41596 27767 41599
rect 28626 41596 28632 41608
rect 27755 41568 28632 41596
rect 27755 41565 27767 41568
rect 27709 41559 27767 41565
rect 28626 41556 28632 41568
rect 28684 41556 28690 41608
rect 28997 41599 29055 41605
rect 28997 41565 29009 41599
rect 29043 41596 29055 41599
rect 29549 41599 29607 41605
rect 29549 41596 29561 41599
rect 29043 41568 29561 41596
rect 29043 41565 29055 41568
rect 28997 41559 29055 41565
rect 29549 41565 29561 41568
rect 29595 41565 29607 41599
rect 29549 41559 29607 41565
rect 29733 41599 29791 41605
rect 29733 41565 29745 41599
rect 29779 41596 29791 41599
rect 30374 41596 30380 41608
rect 29779 41568 30380 41596
rect 29779 41565 29791 41568
rect 29733 41559 29791 41565
rect 30374 41556 30380 41568
rect 30432 41556 30438 41608
rect 30852 41605 30880 41636
rect 31202 41624 31208 41636
rect 31260 41624 31266 41676
rect 37090 41664 37096 41676
rect 37051 41636 37096 41664
rect 37090 41624 37096 41636
rect 37148 41624 37154 41676
rect 30837 41599 30895 41605
rect 30837 41565 30849 41599
rect 30883 41565 30895 41599
rect 30837 41559 30895 41565
rect 31110 41556 31116 41608
rect 31168 41596 31174 41608
rect 31481 41599 31539 41605
rect 31481 41596 31493 41599
rect 31168 41568 31493 41596
rect 31168 41556 31174 41568
rect 31481 41565 31493 41568
rect 31527 41565 31539 41599
rect 31481 41559 31539 41565
rect 34149 41599 34207 41605
rect 34149 41565 34161 41599
rect 34195 41596 34207 41599
rect 34238 41596 34244 41608
rect 34195 41568 34244 41596
rect 34195 41565 34207 41568
rect 34149 41559 34207 41565
rect 34238 41556 34244 41568
rect 34296 41556 34302 41608
rect 34514 41556 34520 41608
rect 34572 41596 34578 41608
rect 36265 41599 36323 41605
rect 36265 41596 36277 41599
rect 34572 41568 36277 41596
rect 34572 41556 34578 41568
rect 36265 41565 36277 41568
rect 36311 41565 36323 41599
rect 36265 41559 36323 41565
rect 21450 41528 21456 41540
rect 20088 41500 21456 41528
rect 21450 41488 21456 41500
rect 21508 41488 21514 41540
rect 30929 41531 30987 41537
rect 30929 41497 30941 41531
rect 30975 41528 30987 41531
rect 31665 41531 31723 41537
rect 31665 41528 31677 41531
rect 30975 41500 31677 41528
rect 30975 41497 30987 41500
rect 30929 41491 30987 41497
rect 31665 41497 31677 41500
rect 31711 41497 31723 41531
rect 31665 41491 31723 41497
rect 33321 41531 33379 41537
rect 33321 41497 33333 41531
rect 33367 41528 33379 41531
rect 34606 41528 34612 41540
rect 33367 41500 34612 41528
rect 33367 41497 33379 41500
rect 33321 41491 33379 41497
rect 34606 41488 34612 41500
rect 34664 41488 34670 41540
rect 36449 41531 36507 41537
rect 36449 41497 36461 41531
rect 36495 41528 36507 41531
rect 37458 41528 37464 41540
rect 36495 41500 37464 41528
rect 36495 41497 36507 41500
rect 36449 41491 36507 41497
rect 37458 41488 37464 41500
rect 37516 41488 37522 41540
rect 17586 41460 17592 41472
rect 10100 41432 17448 41460
rect 17547 41432 17592 41460
rect 10100 41420 10106 41432
rect 17586 41420 17592 41432
rect 17644 41420 17650 41472
rect 17678 41420 17684 41472
rect 17736 41460 17742 41472
rect 20622 41460 20628 41472
rect 17736 41432 20628 41460
rect 17736 41420 17742 41432
rect 20622 41420 20628 41432
rect 20680 41420 20686 41472
rect 26142 41420 26148 41472
rect 26200 41460 26206 41472
rect 26329 41463 26387 41469
rect 26329 41460 26341 41463
rect 26200 41432 26341 41460
rect 26200 41420 26206 41432
rect 26329 41429 26341 41432
rect 26375 41429 26387 41463
rect 26329 41423 26387 41429
rect 28813 41463 28871 41469
rect 28813 41429 28825 41463
rect 28859 41460 28871 41463
rect 28902 41460 28908 41472
rect 28859 41432 28908 41460
rect 28859 41429 28871 41432
rect 28813 41423 28871 41429
rect 28902 41420 28908 41432
rect 28960 41420 28966 41472
rect 1104 41370 38824 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 38824 41370
rect 1104 41296 38824 41318
rect 10502 41256 10508 41268
rect 10463 41228 10508 41256
rect 10502 41216 10508 41228
rect 10560 41256 10566 41268
rect 26878 41256 26884 41268
rect 10560 41228 26884 41256
rect 10560 41216 10566 41228
rect 26878 41216 26884 41228
rect 26936 41216 26942 41268
rect 27157 41259 27215 41265
rect 27157 41225 27169 41259
rect 27203 41256 27215 41259
rect 27706 41256 27712 41268
rect 27203 41228 27712 41256
rect 27203 41225 27215 41228
rect 27157 41219 27215 41225
rect 27706 41216 27712 41228
rect 27764 41216 27770 41268
rect 30006 41256 30012 41268
rect 29967 41228 30012 41256
rect 30006 41216 30012 41228
rect 30064 41216 30070 41268
rect 31110 41256 31116 41268
rect 31071 41228 31116 41256
rect 31110 41216 31116 41228
rect 31168 41216 31174 41268
rect 34238 41256 34244 41268
rect 31726 41228 34100 41256
rect 34199 41228 34244 41256
rect 8757 41191 8815 41197
rect 8757 41157 8769 41191
rect 8803 41188 8815 41191
rect 9217 41191 9275 41197
rect 9217 41188 9229 41191
rect 8803 41160 9229 41188
rect 8803 41157 8815 41160
rect 8757 41151 8815 41157
rect 9217 41157 9229 41160
rect 9263 41188 9275 41191
rect 9674 41188 9680 41200
rect 9263 41160 9680 41188
rect 9263 41157 9275 41160
rect 9217 41151 9275 41157
rect 9674 41148 9680 41160
rect 9732 41148 9738 41200
rect 21266 41148 21272 41200
rect 21324 41188 21330 41200
rect 23382 41188 23388 41200
rect 21324 41160 23388 41188
rect 21324 41148 21330 41160
rect 8386 41120 8392 41132
rect 8347 41092 8392 41120
rect 8386 41080 8392 41092
rect 8444 41080 8450 41132
rect 19426 41120 19432 41132
rect 19387 41092 19432 41120
rect 19426 41080 19432 41092
rect 19484 41080 19490 41132
rect 19705 41123 19763 41129
rect 19705 41089 19717 41123
rect 19751 41120 19763 41123
rect 21174 41120 21180 41132
rect 19751 41092 21180 41120
rect 19751 41089 19763 41092
rect 19705 41083 19763 41089
rect 21174 41080 21180 41092
rect 21232 41080 21238 41132
rect 22664 41129 22692 41160
rect 23382 41148 23388 41160
rect 23440 41148 23446 41200
rect 28902 41197 28908 41200
rect 28896 41188 28908 41197
rect 23952 41160 27108 41188
rect 28863 41160 28908 41188
rect 22649 41123 22707 41129
rect 22649 41089 22661 41123
rect 22695 41089 22707 41123
rect 22649 41083 22707 41089
rect 22738 41080 22744 41132
rect 22796 41120 22802 41132
rect 22905 41123 22963 41129
rect 22905 41120 22917 41123
rect 22796 41092 22917 41120
rect 22796 41080 22802 41092
rect 22905 41089 22917 41092
rect 22951 41089 22963 41123
rect 22905 41083 22963 41089
rect 20622 40876 20628 40928
rect 20680 40916 20686 40928
rect 23952 40916 23980 41160
rect 24949 41123 25007 41129
rect 24949 41089 24961 41123
rect 24995 41120 25007 41123
rect 25222 41120 25228 41132
rect 24995 41092 25228 41120
rect 24995 41089 25007 41092
rect 24949 41083 25007 41089
rect 25222 41080 25228 41092
rect 25280 41080 25286 41132
rect 26970 41120 26976 41132
rect 26931 41092 26976 41120
rect 26970 41080 26976 41092
rect 27028 41080 27034 41132
rect 27080 41120 27108 41160
rect 28896 41151 28908 41160
rect 28902 41148 28908 41151
rect 28960 41148 28966 41200
rect 31726 41188 31754 41228
rect 33042 41188 33048 41200
rect 29012 41160 31754 41188
rect 32416 41160 33048 41188
rect 29012 41120 29040 41160
rect 30926 41120 30932 41132
rect 27080 41092 29040 41120
rect 30887 41092 30932 41120
rect 30926 41080 30932 41092
rect 30984 41080 30990 41132
rect 25133 41055 25191 41061
rect 25133 41021 25145 41055
rect 25179 41021 25191 41055
rect 25133 41015 25191 41021
rect 24029 40987 24087 40993
rect 24029 40953 24041 40987
rect 24075 40984 24087 40987
rect 24854 40984 24860 40996
rect 24075 40956 24860 40984
rect 24075 40953 24087 40956
rect 24029 40947 24087 40953
rect 24854 40944 24860 40956
rect 24912 40984 24918 40996
rect 25148 40984 25176 41015
rect 27982 41012 27988 41064
rect 28040 41052 28046 41064
rect 28626 41052 28632 41064
rect 28040 41024 28632 41052
rect 28040 41012 28046 41024
rect 28626 41012 28632 41024
rect 28684 41012 28690 41064
rect 31754 41012 31760 41064
rect 31812 41052 31818 41064
rect 32416 41061 32444 41160
rect 33042 41148 33048 41160
rect 33100 41148 33106 41200
rect 34072 41188 34100 41228
rect 34238 41216 34244 41228
rect 34296 41216 34302 41268
rect 37458 41256 37464 41268
rect 37419 41228 37464 41256
rect 37458 41216 37464 41228
rect 37516 41216 37522 41268
rect 34072 41160 37412 41188
rect 32674 41129 32680 41132
rect 32668 41083 32680 41129
rect 32732 41120 32738 41132
rect 34425 41123 34483 41129
rect 32732 41092 32768 41120
rect 32674 41080 32680 41083
rect 32732 41080 32738 41092
rect 34425 41089 34437 41123
rect 34471 41120 34483 41123
rect 35253 41123 35311 41129
rect 35253 41120 35265 41123
rect 34471 41092 35265 41120
rect 34471 41089 34483 41092
rect 34425 41083 34483 41089
rect 35253 41089 35265 41092
rect 35299 41120 35311 41123
rect 35986 41120 35992 41132
rect 35299 41092 35992 41120
rect 35299 41089 35311 41092
rect 35253 41083 35311 41089
rect 35986 41080 35992 41092
rect 36044 41080 36050 41132
rect 37384 41129 37412 41160
rect 37369 41123 37427 41129
rect 37369 41089 37381 41123
rect 37415 41089 37427 41123
rect 37369 41083 37427 41089
rect 32401 41055 32459 41061
rect 32401 41052 32413 41055
rect 31812 41024 32413 41052
rect 31812 41012 31818 41024
rect 32401 41021 32413 41024
rect 32447 41021 32459 41055
rect 34609 41055 34667 41061
rect 34609 41052 34621 41055
rect 32401 41015 32459 41021
rect 33796 41024 34621 41052
rect 33796 40993 33824 41024
rect 34609 41021 34621 41024
rect 34655 41052 34667 41055
rect 34790 41052 34796 41064
rect 34655 41024 34796 41052
rect 34655 41021 34667 41024
rect 34609 41015 34667 41021
rect 34790 41012 34796 41024
rect 34848 41012 34854 41064
rect 35069 41055 35127 41061
rect 35069 41021 35081 41055
rect 35115 41052 35127 41055
rect 35342 41052 35348 41064
rect 35115 41024 35348 41052
rect 35115 41021 35127 41024
rect 35069 41015 35127 41021
rect 35342 41012 35348 41024
rect 35400 41012 35406 41064
rect 24912 40956 25176 40984
rect 33781 40987 33839 40993
rect 24912 40944 24918 40956
rect 33781 40953 33793 40987
rect 33827 40953 33839 40987
rect 38378 40984 38384 40996
rect 33781 40947 33839 40953
rect 35360 40956 38384 40984
rect 20680 40888 23980 40916
rect 24765 40919 24823 40925
rect 20680 40876 20686 40888
rect 24765 40885 24777 40919
rect 24811 40916 24823 40919
rect 25130 40916 25136 40928
rect 24811 40888 25136 40916
rect 24811 40885 24823 40888
rect 24765 40879 24823 40885
rect 25130 40876 25136 40888
rect 25188 40876 25194 40928
rect 26878 40876 26884 40928
rect 26936 40916 26942 40928
rect 35360 40916 35388 40956
rect 38378 40944 38384 40956
rect 38436 40944 38442 40996
rect 26936 40888 35388 40916
rect 35437 40919 35495 40925
rect 26936 40876 26942 40888
rect 35437 40885 35449 40919
rect 35483 40916 35495 40919
rect 35802 40916 35808 40928
rect 35483 40888 35808 40916
rect 35483 40885 35495 40888
rect 35437 40879 35495 40885
rect 35802 40876 35808 40888
rect 35860 40876 35866 40928
rect 36078 40916 36084 40928
rect 36039 40888 36084 40916
rect 36078 40876 36084 40888
rect 36136 40876 36142 40928
rect 36262 40876 36268 40928
rect 36320 40916 36326 40928
rect 36541 40919 36599 40925
rect 36541 40916 36553 40919
rect 36320 40888 36553 40916
rect 36320 40876 36326 40888
rect 36541 40885 36553 40888
rect 36587 40885 36599 40919
rect 36541 40879 36599 40885
rect 1104 40826 38824 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 38824 40826
rect 1104 40752 38824 40774
rect 20993 40715 21051 40721
rect 20993 40681 21005 40715
rect 21039 40712 21051 40715
rect 21266 40712 21272 40724
rect 21039 40684 21272 40712
rect 21039 40681 21051 40684
rect 20993 40675 21051 40681
rect 21266 40672 21272 40684
rect 21324 40672 21330 40724
rect 23477 40715 23535 40721
rect 23477 40681 23489 40715
rect 23523 40712 23535 40715
rect 23658 40712 23664 40724
rect 23523 40684 23664 40712
rect 23523 40681 23535 40684
rect 23477 40675 23535 40681
rect 23658 40672 23664 40684
rect 23716 40672 23722 40724
rect 25133 40715 25191 40721
rect 25133 40681 25145 40715
rect 25179 40712 25191 40715
rect 26050 40712 26056 40724
rect 25179 40684 26056 40712
rect 25179 40681 25191 40684
rect 25133 40675 25191 40681
rect 26050 40672 26056 40684
rect 26108 40672 26114 40724
rect 32674 40712 32680 40724
rect 32635 40684 32680 40712
rect 32674 40672 32680 40684
rect 32732 40672 32738 40724
rect 34149 40715 34207 40721
rect 34149 40681 34161 40715
rect 34195 40712 34207 40715
rect 34514 40712 34520 40724
rect 34195 40684 34520 40712
rect 34195 40681 34207 40684
rect 34149 40675 34207 40681
rect 34514 40672 34520 40684
rect 34572 40672 34578 40724
rect 34698 40672 34704 40724
rect 34756 40712 34762 40724
rect 34885 40715 34943 40721
rect 34885 40712 34897 40715
rect 34756 40684 34897 40712
rect 34756 40672 34762 40684
rect 34885 40681 34897 40684
rect 34931 40681 34943 40715
rect 34885 40675 34943 40681
rect 10962 40536 10968 40588
rect 11020 40576 11026 40588
rect 11425 40579 11483 40585
rect 11425 40576 11437 40579
rect 11020 40548 11437 40576
rect 11020 40536 11026 40548
rect 11425 40545 11437 40548
rect 11471 40576 11483 40579
rect 15286 40576 15292 40588
rect 11471 40548 15292 40576
rect 11471 40545 11483 40548
rect 11425 40539 11483 40545
rect 15286 40536 15292 40548
rect 15344 40536 15350 40588
rect 18690 40536 18696 40588
rect 18748 40576 18754 40588
rect 19521 40579 19579 40585
rect 19521 40576 19533 40579
rect 18748 40548 19533 40576
rect 18748 40536 18754 40548
rect 19521 40545 19533 40548
rect 19567 40545 19579 40579
rect 21284 40576 21312 40672
rect 25777 40647 25835 40653
rect 25777 40613 25789 40647
rect 25823 40644 25835 40647
rect 25866 40644 25872 40656
rect 25823 40616 25872 40644
rect 25823 40613 25835 40616
rect 25777 40607 25835 40613
rect 21637 40579 21695 40585
rect 21637 40576 21649 40579
rect 21284 40548 21649 40576
rect 19521 40539 19579 40545
rect 21637 40545 21649 40548
rect 21683 40545 21695 40579
rect 21637 40539 21695 40545
rect 24765 40579 24823 40585
rect 24765 40545 24777 40579
rect 24811 40576 24823 40579
rect 24854 40576 24860 40588
rect 24811 40548 24860 40576
rect 24811 40545 24823 40548
rect 24765 40539 24823 40545
rect 24854 40536 24860 40548
rect 24912 40536 24918 40588
rect 24974 40579 25032 40585
rect 24974 40545 24986 40579
rect 25020 40576 25032 40579
rect 25792 40576 25820 40607
rect 25866 40604 25872 40616
rect 25924 40644 25930 40656
rect 26142 40644 26148 40656
rect 25924 40616 26148 40644
rect 25924 40604 25930 40616
rect 26142 40604 26148 40616
rect 26200 40604 26206 40656
rect 25020 40548 25820 40576
rect 25020 40545 25032 40548
rect 24974 40539 25032 40545
rect 34606 40536 34612 40588
rect 34664 40576 34670 40588
rect 34977 40579 35035 40585
rect 34977 40576 34989 40579
rect 34664 40548 34989 40576
rect 34664 40536 34670 40548
rect 34977 40545 34989 40548
rect 35023 40545 35035 40579
rect 36262 40576 36268 40588
rect 36223 40548 36268 40576
rect 34977 40539 35035 40545
rect 36262 40536 36268 40548
rect 36320 40536 36326 40588
rect 38105 40579 38163 40585
rect 38105 40545 38117 40579
rect 38151 40576 38163 40579
rect 38194 40576 38200 40588
rect 38151 40548 38200 40576
rect 38151 40545 38163 40548
rect 38105 40539 38163 40545
rect 38194 40536 38200 40548
rect 38252 40536 38258 40588
rect 1578 40508 1584 40520
rect 1539 40480 1584 40508
rect 1578 40468 1584 40480
rect 1636 40468 1642 40520
rect 9674 40508 9680 40520
rect 9635 40480 9680 40508
rect 9674 40468 9680 40480
rect 9732 40468 9738 40520
rect 16485 40511 16543 40517
rect 16485 40477 16497 40511
rect 16531 40508 16543 40511
rect 16758 40508 16764 40520
rect 16531 40480 16764 40508
rect 16531 40477 16543 40480
rect 16485 40471 16543 40477
rect 16758 40468 16764 40480
rect 16816 40468 16822 40520
rect 19245 40511 19303 40517
rect 19245 40477 19257 40511
rect 19291 40508 19303 40511
rect 21174 40508 21180 40520
rect 19291 40480 21180 40508
rect 19291 40477 19303 40480
rect 19245 40471 19303 40477
rect 21174 40468 21180 40480
rect 21232 40468 21238 40520
rect 23658 40508 23664 40520
rect 23619 40480 23664 40508
rect 23658 40468 23664 40480
rect 23716 40468 23722 40520
rect 23845 40511 23903 40517
rect 23845 40477 23857 40511
rect 23891 40508 23903 40511
rect 24489 40511 24547 40517
rect 24489 40508 24501 40511
rect 23891 40480 24501 40508
rect 23891 40477 23903 40480
rect 23845 40471 23903 40477
rect 24489 40477 24501 40480
rect 24535 40508 24547 40511
rect 26053 40511 26111 40517
rect 26053 40508 26065 40511
rect 24535 40480 26065 40508
rect 24535 40477 24547 40480
rect 24489 40471 24547 40477
rect 21082 40440 21088 40452
rect 21043 40412 21088 40440
rect 21082 40400 21088 40412
rect 21140 40400 21146 40452
rect 21904 40443 21962 40449
rect 21904 40409 21916 40443
rect 21950 40440 21962 40443
rect 22094 40440 22100 40452
rect 21950 40412 22100 40440
rect 21950 40409 21962 40412
rect 21904 40403 21962 40409
rect 22094 40400 22100 40412
rect 22152 40400 22158 40452
rect 16666 40372 16672 40384
rect 16627 40344 16672 40372
rect 16666 40332 16672 40344
rect 16724 40332 16730 40384
rect 23017 40375 23075 40381
rect 23017 40341 23029 40375
rect 23063 40372 23075 40375
rect 23860 40372 23888 40471
rect 24964 40452 24992 40480
rect 26053 40477 26065 40480
rect 26099 40477 26111 40511
rect 26053 40471 26111 40477
rect 27706 40468 27712 40520
rect 27764 40517 27770 40520
rect 27764 40508 27776 40517
rect 27982 40508 27988 40520
rect 27764 40480 27809 40508
rect 27943 40480 27988 40508
rect 27764 40471 27776 40480
rect 27764 40468 27770 40471
rect 27982 40468 27988 40480
rect 28040 40468 28046 40520
rect 32858 40508 32864 40520
rect 32819 40480 32864 40508
rect 32858 40468 32864 40480
rect 32916 40468 32922 40520
rect 34790 40468 34796 40520
rect 34848 40508 34854 40520
rect 34885 40511 34943 40517
rect 34885 40508 34897 40511
rect 34848 40480 34897 40508
rect 34848 40468 34854 40480
rect 34885 40477 34897 40480
rect 34931 40477 34943 40511
rect 35802 40508 35808 40520
rect 35763 40480 35808 40508
rect 34885 40471 34943 40477
rect 35802 40468 35808 40480
rect 35860 40468 35866 40520
rect 24946 40400 24952 40452
rect 25004 40400 25010 40452
rect 25222 40440 25228 40452
rect 25056 40412 25228 40440
rect 23063 40344 23888 40372
rect 24857 40375 24915 40381
rect 23063 40341 23075 40344
rect 23017 40335 23075 40341
rect 24857 40341 24869 40375
rect 24903 40372 24915 40375
rect 25056 40372 25084 40412
rect 25222 40400 25228 40412
rect 25280 40440 25286 40452
rect 35161 40443 35219 40449
rect 25280 40412 25820 40440
rect 25280 40400 25286 40412
rect 25792 40384 25820 40412
rect 35161 40409 35173 40443
rect 35207 40440 35219 40443
rect 35342 40440 35348 40452
rect 35207 40412 35348 40440
rect 35207 40409 35219 40412
rect 35161 40403 35219 40409
rect 35342 40400 35348 40412
rect 35400 40400 35406 40452
rect 36449 40443 36507 40449
rect 36449 40409 36461 40443
rect 36495 40440 36507 40443
rect 37366 40440 37372 40452
rect 36495 40412 37372 40440
rect 36495 40409 36507 40412
rect 36449 40403 36507 40409
rect 37366 40400 37372 40412
rect 37424 40400 37430 40452
rect 25590 40372 25596 40384
rect 24903 40344 25084 40372
rect 25551 40344 25596 40372
rect 24903 40341 24915 40344
rect 24857 40335 24915 40341
rect 25590 40332 25596 40344
rect 25648 40332 25654 40384
rect 25774 40332 25780 40384
rect 25832 40372 25838 40384
rect 26605 40375 26663 40381
rect 26605 40372 26617 40375
rect 25832 40344 26617 40372
rect 25832 40332 25838 40344
rect 26605 40341 26617 40344
rect 26651 40341 26663 40375
rect 26605 40335 26663 40341
rect 33594 40332 33600 40384
rect 33652 40372 33658 40384
rect 34701 40375 34759 40381
rect 34701 40372 34713 40375
rect 33652 40344 34713 40372
rect 33652 40332 33658 40344
rect 34701 40341 34713 40344
rect 34747 40341 34759 40375
rect 35618 40372 35624 40384
rect 35579 40344 35624 40372
rect 34701 40335 34759 40341
rect 35618 40332 35624 40344
rect 35676 40332 35682 40384
rect 1104 40282 38824 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 38824 40282
rect 1104 40208 38824 40230
rect 9766 40128 9772 40180
rect 9824 40168 9830 40180
rect 9824 40140 17816 40168
rect 9824 40128 9830 40140
rect 3418 40100 3424 40112
rect 3379 40072 3424 40100
rect 3418 40060 3424 40072
rect 3476 40060 3482 40112
rect 9674 40060 9680 40112
rect 9732 40100 9738 40112
rect 10520 40109 10548 40140
rect 10505 40103 10563 40109
rect 9732 40072 9812 40100
rect 9732 40060 9738 40072
rect 1578 40032 1584 40044
rect 1539 40004 1584 40032
rect 1578 39992 1584 40004
rect 1636 39992 1642 40044
rect 9784 40041 9812 40072
rect 10505 40069 10517 40103
rect 10551 40069 10563 40103
rect 10505 40063 10563 40069
rect 16666 40060 16672 40112
rect 16724 40100 16730 40112
rect 16914 40103 16972 40109
rect 16914 40100 16926 40103
rect 16724 40072 16926 40100
rect 16724 40060 16730 40072
rect 16914 40069 16926 40072
rect 16960 40069 16972 40103
rect 17788 40100 17816 40140
rect 17862 40128 17868 40180
rect 17920 40168 17926 40180
rect 18049 40171 18107 40177
rect 18049 40168 18061 40171
rect 17920 40140 18061 40168
rect 17920 40128 17926 40140
rect 18049 40137 18061 40140
rect 18095 40137 18107 40171
rect 18049 40131 18107 40137
rect 19889 40171 19947 40177
rect 19889 40137 19901 40171
rect 19935 40168 19947 40171
rect 20346 40168 20352 40180
rect 19935 40140 20352 40168
rect 19935 40137 19947 40140
rect 19889 40131 19947 40137
rect 20346 40128 20352 40140
rect 20404 40128 20410 40180
rect 23658 40128 23664 40180
rect 23716 40168 23722 40180
rect 23716 40140 26004 40168
rect 23716 40128 23722 40140
rect 22646 40100 22652 40112
rect 17788 40072 22652 40100
rect 16914 40063 16972 40069
rect 22646 40060 22652 40072
rect 22704 40060 22710 40112
rect 25133 40103 25191 40109
rect 25133 40069 25145 40103
rect 25179 40100 25191 40103
rect 25976 40100 26004 40140
rect 26970 40128 26976 40180
rect 27028 40168 27034 40180
rect 27341 40171 27399 40177
rect 27341 40168 27353 40171
rect 27028 40140 27353 40168
rect 27028 40128 27034 40140
rect 27341 40137 27353 40140
rect 27387 40137 27399 40171
rect 27341 40131 27399 40137
rect 30193 40171 30251 40177
rect 30193 40137 30205 40171
rect 30239 40168 30251 40171
rect 30650 40168 30656 40180
rect 30239 40140 30656 40168
rect 30239 40137 30251 40140
rect 30193 40131 30251 40137
rect 30650 40128 30656 40140
rect 30708 40128 30714 40180
rect 30742 40100 30748 40112
rect 25179 40072 25912 40100
rect 25976 40072 27200 40100
rect 30703 40072 30748 40100
rect 25179 40069 25191 40072
rect 25133 40063 25191 40069
rect 25884 40044 25912 40072
rect 9769 40035 9827 40041
rect 9769 40001 9781 40035
rect 9815 40001 9827 40035
rect 9769 39995 9827 40001
rect 18138 39992 18144 40044
rect 18196 40032 18202 40044
rect 18765 40035 18823 40041
rect 18765 40032 18777 40035
rect 18196 40004 18777 40032
rect 18196 39992 18202 40004
rect 18765 40001 18777 40004
rect 18811 40001 18823 40035
rect 20346 40032 20352 40044
rect 20307 40004 20352 40032
rect 18765 39995 18823 40001
rect 20346 39992 20352 40004
rect 20404 39992 20410 40044
rect 20533 40035 20591 40041
rect 20533 40001 20545 40035
rect 20579 40001 20591 40035
rect 20533 39995 20591 40001
rect 1762 39964 1768 39976
rect 1723 39936 1768 39964
rect 1762 39924 1768 39936
rect 1820 39924 1826 39976
rect 16669 39967 16727 39973
rect 16669 39933 16681 39967
rect 16715 39933 16727 39967
rect 16669 39927 16727 39933
rect 18509 39967 18567 39973
rect 18509 39933 18521 39967
rect 18555 39933 18567 39967
rect 18509 39927 18567 39933
rect 16684 39828 16712 39927
rect 18524 39828 18552 39927
rect 19518 39924 19524 39976
rect 19576 39964 19582 39976
rect 20548 39964 20576 39995
rect 21174 39992 21180 40044
rect 21232 40032 21238 40044
rect 21910 40032 21916 40044
rect 21232 40004 21916 40032
rect 21232 39992 21238 40004
rect 21910 39992 21916 40004
rect 21968 40032 21974 40044
rect 22097 40035 22155 40041
rect 22097 40032 22109 40035
rect 21968 40004 22109 40032
rect 21968 39992 21974 40004
rect 22097 40001 22109 40004
rect 22143 40001 22155 40035
rect 22097 39995 22155 40001
rect 24854 39992 24860 40044
rect 24912 40032 24918 40044
rect 25593 40035 25651 40041
rect 25593 40032 25605 40035
rect 24912 40004 25605 40032
rect 24912 39992 24918 40004
rect 25593 40001 25605 40004
rect 25639 40001 25651 40035
rect 25774 40032 25780 40044
rect 25735 40004 25780 40032
rect 25593 39995 25651 40001
rect 25774 39992 25780 40004
rect 25832 39992 25838 40044
rect 25866 39992 25872 40044
rect 25924 40032 25930 40044
rect 27172 40041 27200 40072
rect 30742 40060 30748 40072
rect 30800 40060 30806 40112
rect 26973 40035 27031 40041
rect 26973 40032 26985 40035
rect 25924 40004 26985 40032
rect 25924 39992 25930 40004
rect 26973 40001 26985 40004
rect 27019 40001 27031 40035
rect 26973 39995 27031 40001
rect 27157 40035 27215 40041
rect 27157 40001 27169 40035
rect 27203 40001 27215 40035
rect 27157 39995 27215 40001
rect 27982 39992 27988 40044
rect 28040 40032 28046 40044
rect 28813 40035 28871 40041
rect 28813 40032 28825 40035
rect 28040 40004 28825 40032
rect 28040 39992 28046 40004
rect 28813 40001 28825 40004
rect 28859 40001 28871 40035
rect 28813 39995 28871 40001
rect 20622 39964 20628 39976
rect 19576 39936 20628 39964
rect 19576 39924 19582 39936
rect 20622 39924 20628 39936
rect 20680 39924 20686 39976
rect 20990 39924 20996 39976
rect 21048 39964 21054 39976
rect 21821 39967 21879 39973
rect 21821 39964 21833 39967
rect 21048 39936 21833 39964
rect 21048 39924 21054 39936
rect 21821 39933 21833 39936
rect 21867 39964 21879 39967
rect 23658 39964 23664 39976
rect 21867 39936 23664 39964
rect 21867 39933 21879 39936
rect 21821 39927 21879 39933
rect 23658 39924 23664 39936
rect 23716 39924 23722 39976
rect 21266 39896 21272 39908
rect 19444 39868 21272 39896
rect 19444 39828 19472 39868
rect 21266 39856 21272 39868
rect 21324 39856 21330 39908
rect 24857 39899 24915 39905
rect 24857 39865 24869 39899
rect 24903 39896 24915 39899
rect 24946 39896 24952 39908
rect 24903 39868 24952 39896
rect 24903 39865 24915 39868
rect 24857 39859 24915 39865
rect 24946 39856 24952 39868
rect 25004 39856 25010 39908
rect 16684 39800 19472 39828
rect 20717 39831 20775 39837
rect 20717 39797 20729 39831
rect 20763 39828 20775 39831
rect 20806 39828 20812 39840
rect 20763 39800 20812 39828
rect 20763 39797 20775 39800
rect 20717 39791 20775 39797
rect 20806 39788 20812 39800
rect 20864 39788 20870 39840
rect 24670 39828 24676 39840
rect 24631 39800 24676 39828
rect 24670 39788 24676 39800
rect 24728 39788 24734 39840
rect 25774 39828 25780 39840
rect 25735 39800 25780 39828
rect 25774 39788 25780 39800
rect 25832 39788 25838 39840
rect 28828 39828 28856 39995
rect 28902 39992 28908 40044
rect 28960 40032 28966 40044
rect 29069 40035 29127 40041
rect 29069 40032 29081 40035
rect 28960 40004 29081 40032
rect 28960 39992 28966 40004
rect 29069 40001 29081 40004
rect 29115 40001 29127 40035
rect 31570 40032 31576 40044
rect 31531 40004 31576 40032
rect 29069 39995 29127 40001
rect 31570 39992 31576 40004
rect 31628 39992 31634 40044
rect 31754 40032 31760 40044
rect 31726 39992 31760 40032
rect 31812 39992 31818 40044
rect 33226 40032 33232 40044
rect 33284 40041 33290 40044
rect 34238 40041 34244 40044
rect 33196 40004 33232 40032
rect 33226 39992 33232 40004
rect 33284 39995 33296 40041
rect 34232 39995 34244 40041
rect 34296 40032 34302 40044
rect 34296 40004 34332 40032
rect 33284 39992 33290 39995
rect 34238 39992 34244 39995
rect 34296 39992 34302 40004
rect 34698 39992 34704 40044
rect 34756 40032 34762 40044
rect 35986 40032 35992 40044
rect 34756 40004 35848 40032
rect 35947 40004 35992 40032
rect 34756 39992 34762 40004
rect 30929 39899 30987 39905
rect 30929 39896 30941 39899
rect 29748 39868 30941 39896
rect 29748 39828 29776 39868
rect 30929 39865 30941 39868
rect 30975 39896 30987 39899
rect 31726 39896 31754 39992
rect 33505 39967 33563 39973
rect 33505 39933 33517 39967
rect 33551 39964 33563 39967
rect 33962 39964 33968 39976
rect 33551 39936 33968 39964
rect 33551 39933 33563 39936
rect 33505 39927 33563 39933
rect 33962 39924 33968 39936
rect 34020 39924 34026 39976
rect 35820 39964 35848 40004
rect 35986 39992 35992 40004
rect 36044 39992 36050 40044
rect 37277 40035 37335 40041
rect 37277 40001 37289 40035
rect 37323 40001 37335 40035
rect 37277 39995 37335 40001
rect 36173 39967 36231 39973
rect 36173 39964 36185 39967
rect 35820 39936 36185 39964
rect 36173 39933 36185 39936
rect 36219 39933 36231 39967
rect 37292 39964 37320 39995
rect 37366 39992 37372 40044
rect 37424 40032 37430 40044
rect 37424 40004 37469 40032
rect 37424 39992 37430 40004
rect 37918 39964 37924 39976
rect 37292 39936 37924 39964
rect 36173 39927 36231 39933
rect 37918 39924 37924 39936
rect 37976 39924 37982 39976
rect 30975 39868 31754 39896
rect 30975 39865 30987 39868
rect 30929 39859 30987 39865
rect 31386 39828 31392 39840
rect 28828 39800 29776 39828
rect 31347 39800 31392 39828
rect 31386 39788 31392 39800
rect 31444 39788 31450 39840
rect 32122 39828 32128 39840
rect 32083 39800 32128 39828
rect 32122 39788 32128 39800
rect 32180 39788 32186 39840
rect 35342 39828 35348 39840
rect 35303 39800 35348 39828
rect 35342 39788 35348 39800
rect 35400 39788 35406 39840
rect 35802 39828 35808 39840
rect 35763 39800 35808 39828
rect 35802 39788 35808 39800
rect 35860 39788 35866 39840
rect 38105 39831 38163 39837
rect 38105 39797 38117 39831
rect 38151 39828 38163 39831
rect 38194 39828 38200 39840
rect 38151 39800 38200 39828
rect 38151 39797 38163 39800
rect 38105 39791 38163 39797
rect 38194 39788 38200 39800
rect 38252 39788 38258 39840
rect 1104 39738 38824 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 38824 39738
rect 1104 39664 38824 39686
rect 1762 39584 1768 39636
rect 1820 39624 1826 39636
rect 2041 39627 2099 39633
rect 2041 39624 2053 39627
rect 1820 39596 2053 39624
rect 1820 39584 1826 39596
rect 2041 39593 2053 39596
rect 2087 39593 2099 39627
rect 16758 39624 16764 39636
rect 16719 39596 16764 39624
rect 2041 39587 2099 39593
rect 16758 39584 16764 39596
rect 16816 39584 16822 39636
rect 18138 39624 18144 39636
rect 18099 39596 18144 39624
rect 18138 39584 18144 39596
rect 18196 39584 18202 39636
rect 24857 39627 24915 39633
rect 24857 39593 24869 39627
rect 24903 39624 24915 39627
rect 25038 39624 25044 39636
rect 24903 39596 25044 39624
rect 24903 39593 24915 39596
rect 24857 39587 24915 39593
rect 25038 39584 25044 39596
rect 25096 39624 25102 39636
rect 25590 39624 25596 39636
rect 25096 39596 25596 39624
rect 25096 39584 25102 39596
rect 25590 39584 25596 39596
rect 25648 39584 25654 39636
rect 28537 39627 28595 39633
rect 28537 39593 28549 39627
rect 28583 39624 28595 39627
rect 28902 39624 28908 39636
rect 28583 39596 28908 39624
rect 28583 39593 28595 39596
rect 28537 39587 28595 39593
rect 28902 39584 28908 39596
rect 28960 39584 28966 39636
rect 31113 39627 31171 39633
rect 31113 39593 31125 39627
rect 31159 39624 31171 39627
rect 31570 39624 31576 39636
rect 31159 39596 31576 39624
rect 31159 39593 31171 39596
rect 31113 39587 31171 39593
rect 31570 39584 31576 39596
rect 31628 39584 31634 39636
rect 32401 39627 32459 39633
rect 32401 39593 32413 39627
rect 32447 39624 32459 39627
rect 32858 39624 32864 39636
rect 32447 39596 32864 39624
rect 32447 39593 32459 39596
rect 32401 39587 32459 39593
rect 32858 39584 32864 39596
rect 32916 39584 32922 39636
rect 33045 39627 33103 39633
rect 33045 39593 33057 39627
rect 33091 39624 33103 39627
rect 33226 39624 33232 39636
rect 33091 39596 33232 39624
rect 33091 39593 33103 39596
rect 33045 39587 33103 39593
rect 33226 39584 33232 39596
rect 33284 39584 33290 39636
rect 34149 39627 34207 39633
rect 34149 39593 34161 39627
rect 34195 39624 34207 39627
rect 34238 39624 34244 39636
rect 34195 39596 34244 39624
rect 34195 39593 34207 39596
rect 34149 39587 34207 39593
rect 34238 39584 34244 39596
rect 34296 39584 34302 39636
rect 35802 39624 35808 39636
rect 34624 39596 35808 39624
rect 17129 39491 17187 39497
rect 17129 39457 17141 39491
rect 17175 39488 17187 39491
rect 17586 39488 17592 39500
rect 17175 39460 17592 39488
rect 17175 39457 17187 39460
rect 17129 39451 17187 39457
rect 17586 39448 17592 39460
rect 17644 39448 17650 39500
rect 21177 39491 21235 39497
rect 21177 39457 21189 39491
rect 21223 39488 21235 39491
rect 21266 39488 21272 39500
rect 21223 39460 21272 39488
rect 21223 39457 21235 39460
rect 21177 39451 21235 39457
rect 21266 39448 21272 39460
rect 21324 39448 21330 39500
rect 25774 39488 25780 39500
rect 21836 39460 22094 39488
rect 2130 39420 2136 39432
rect 2091 39392 2136 39420
rect 2130 39380 2136 39392
rect 2188 39380 2194 39432
rect 16945 39423 17003 39429
rect 16945 39389 16957 39423
rect 16991 39389 17003 39423
rect 16945 39383 17003 39389
rect 17957 39423 18015 39429
rect 17957 39389 17969 39423
rect 18003 39420 18015 39423
rect 18322 39420 18328 39432
rect 18003 39392 18328 39420
rect 18003 39389 18015 39392
rect 17957 39383 18015 39389
rect 16850 39312 16856 39364
rect 16908 39352 16914 39364
rect 16960 39352 16988 39383
rect 18322 39380 18328 39392
rect 18380 39380 18386 39432
rect 18690 39352 18696 39364
rect 16908 39324 18696 39352
rect 16908 39312 16914 39324
rect 18690 39312 18696 39324
rect 18748 39312 18754 39364
rect 20898 39352 20904 39364
rect 20956 39361 20962 39364
rect 20868 39324 20904 39352
rect 20898 39312 20904 39324
rect 20956 39315 20968 39361
rect 20956 39312 20962 39315
rect 21836 39296 21864 39460
rect 21910 39380 21916 39432
rect 21968 39420 21974 39432
rect 21968 39392 22013 39420
rect 21968 39380 21974 39392
rect 22066 39352 22094 39460
rect 25056 39460 25780 39488
rect 24670 39380 24676 39432
rect 24728 39420 24734 39432
rect 25056 39429 25084 39460
rect 25774 39448 25780 39460
rect 25832 39448 25838 39500
rect 30650 39448 30656 39500
rect 30708 39488 30714 39500
rect 30745 39491 30803 39497
rect 30745 39488 30757 39491
rect 30708 39460 30757 39488
rect 30708 39448 30714 39460
rect 30745 39457 30757 39460
rect 30791 39457 30803 39491
rect 30745 39451 30803 39457
rect 24765 39423 24823 39429
rect 24765 39420 24777 39423
rect 24728 39392 24777 39420
rect 24728 39380 24734 39392
rect 24765 39389 24777 39392
rect 24811 39389 24823 39423
rect 24765 39383 24823 39389
rect 25041 39423 25099 39429
rect 25041 39389 25053 39423
rect 25087 39389 25099 39423
rect 25041 39383 25099 39389
rect 25130 39380 25136 39432
rect 25188 39420 25194 39432
rect 28350 39420 28356 39432
rect 25188 39392 25233 39420
rect 28311 39392 28356 39420
rect 25188 39380 25194 39392
rect 28350 39380 28356 39392
rect 28408 39380 28414 39432
rect 30929 39423 30987 39429
rect 30929 39389 30941 39423
rect 30975 39420 30987 39423
rect 32122 39420 32128 39432
rect 30975 39392 31754 39420
rect 32083 39392 32128 39420
rect 30975 39389 30987 39392
rect 30929 39383 30987 39389
rect 29546 39352 29552 39364
rect 22066 39324 29552 39352
rect 29546 39312 29552 39324
rect 29604 39312 29610 39364
rect 31726 39352 31754 39392
rect 32122 39380 32128 39392
rect 32180 39380 32186 39432
rect 32217 39423 32275 39429
rect 32217 39389 32229 39423
rect 32263 39420 32275 39423
rect 32306 39420 32312 39432
rect 32263 39392 32312 39420
rect 32263 39389 32275 39392
rect 32217 39383 32275 39389
rect 32232 39352 32260 39383
rect 32306 39380 32312 39392
rect 32364 39380 32370 39432
rect 32490 39380 32496 39432
rect 32548 39420 32554 39432
rect 32861 39423 32919 39429
rect 32861 39420 32873 39423
rect 32548 39392 32873 39420
rect 32548 39380 32554 39392
rect 32861 39389 32873 39392
rect 32907 39389 32919 39423
rect 32861 39383 32919 39389
rect 33965 39423 34023 39429
rect 33965 39389 33977 39423
rect 34011 39420 34023 39423
rect 34624 39420 34652 39596
rect 35802 39584 35808 39596
rect 35860 39584 35866 39636
rect 34790 39516 34796 39568
rect 34848 39556 34854 39568
rect 35253 39559 35311 39565
rect 35253 39556 35265 39559
rect 34848 39528 35265 39556
rect 34848 39516 34854 39528
rect 35253 39525 35265 39528
rect 35299 39525 35311 39559
rect 35253 39519 35311 39525
rect 34698 39448 34704 39500
rect 34756 39488 34762 39500
rect 34756 39460 35112 39488
rect 34756 39448 34762 39460
rect 35084 39429 35112 39460
rect 36078 39448 36084 39500
rect 36136 39488 36142 39500
rect 36265 39491 36323 39497
rect 36265 39488 36277 39491
rect 36136 39460 36277 39488
rect 36136 39448 36142 39460
rect 36265 39457 36277 39460
rect 36311 39457 36323 39491
rect 38102 39488 38108 39500
rect 38063 39460 38108 39488
rect 36265 39451 36323 39457
rect 38102 39448 38108 39460
rect 38160 39448 38166 39500
rect 34011 39392 34652 39420
rect 35069 39423 35127 39429
rect 34011 39389 34023 39392
rect 33965 39383 34023 39389
rect 35069 39389 35081 39423
rect 35115 39389 35127 39423
rect 35069 39383 35127 39389
rect 31726 39324 32260 39352
rect 34606 39312 34612 39364
rect 34664 39352 34670 39364
rect 34885 39355 34943 39361
rect 34664 39324 34836 39352
rect 34664 39312 34670 39324
rect 19797 39287 19855 39293
rect 19797 39253 19809 39287
rect 19843 39284 19855 39287
rect 20070 39284 20076 39296
rect 19843 39256 20076 39284
rect 19843 39253 19855 39256
rect 19797 39247 19855 39253
rect 20070 39244 20076 39256
rect 20128 39244 20134 39296
rect 21729 39287 21787 39293
rect 21729 39253 21741 39287
rect 21775 39284 21787 39287
rect 21818 39284 21824 39296
rect 21775 39256 21824 39284
rect 21775 39253 21787 39256
rect 21729 39247 21787 39253
rect 21818 39244 21824 39256
rect 21876 39244 21882 39296
rect 25314 39284 25320 39296
rect 25275 39256 25320 39284
rect 25314 39244 25320 39256
rect 25372 39244 25378 39296
rect 34698 39284 34704 39296
rect 34659 39256 34704 39284
rect 34698 39244 34704 39256
rect 34756 39244 34762 39296
rect 34808 39284 34836 39324
rect 34885 39321 34897 39355
rect 34931 39352 34943 39355
rect 36446 39352 36452 39364
rect 34931 39324 35204 39352
rect 36407 39324 36452 39352
rect 34931 39321 34943 39324
rect 34885 39315 34943 39321
rect 34974 39284 34980 39296
rect 34808 39256 34980 39284
rect 34974 39244 34980 39256
rect 35032 39244 35038 39296
rect 35176 39284 35204 39324
rect 36446 39312 36452 39324
rect 36504 39312 36510 39364
rect 35342 39284 35348 39296
rect 35176 39256 35348 39284
rect 35342 39244 35348 39256
rect 35400 39244 35406 39296
rect 1104 39194 38824 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 38824 39194
rect 1104 39120 38824 39142
rect 18322 39080 18328 39092
rect 18283 39052 18328 39080
rect 18322 39040 18328 39052
rect 18380 39040 18386 39092
rect 20898 39040 20904 39092
rect 20956 39080 20962 39092
rect 20993 39083 21051 39089
rect 20993 39080 21005 39083
rect 20956 39052 21005 39080
rect 20956 39040 20962 39052
rect 20993 39049 21005 39052
rect 21039 39049 21051 39083
rect 20993 39043 21051 39049
rect 22189 39083 22247 39089
rect 22189 39049 22201 39083
rect 22235 39080 22247 39083
rect 28350 39080 28356 39092
rect 22235 39052 28356 39080
rect 22235 39049 22247 39052
rect 22189 39043 22247 39049
rect 28350 39040 28356 39052
rect 28408 39040 28414 39092
rect 32490 39080 32496 39092
rect 32451 39052 32496 39080
rect 32490 39040 32496 39052
rect 32548 39040 32554 39092
rect 36446 39040 36452 39092
rect 36504 39080 36510 39092
rect 37553 39083 37611 39089
rect 37553 39080 37565 39083
rect 36504 39052 37565 39080
rect 36504 39040 36510 39052
rect 37553 39049 37565 39052
rect 37599 39049 37611 39083
rect 37553 39043 37611 39049
rect 1670 38972 1676 39024
rect 1728 39012 1734 39024
rect 19426 39012 19432 39024
rect 1728 38984 6914 39012
rect 1728 38972 1734 38984
rect 6886 38944 6914 38984
rect 18524 38984 19432 39012
rect 14277 38947 14335 38953
rect 14277 38944 14289 38947
rect 6886 38916 14289 38944
rect 14277 38913 14289 38916
rect 14323 38913 14335 38947
rect 16850 38944 16856 38956
rect 16811 38916 16856 38944
rect 14277 38907 14335 38913
rect 16850 38904 16856 38916
rect 16908 38904 16914 38956
rect 18524 38953 18552 38984
rect 19426 38972 19432 38984
rect 19484 38972 19490 39024
rect 25869 39015 25927 39021
rect 25869 39012 25881 39015
rect 24780 38984 25881 39012
rect 18509 38947 18567 38953
rect 18509 38913 18521 38947
rect 18555 38913 18567 38947
rect 18509 38907 18567 38913
rect 18598 38904 18604 38956
rect 18656 38944 18662 38956
rect 19978 38944 19984 38956
rect 18656 38916 18701 38944
rect 19939 38916 19984 38944
rect 18656 38904 18662 38916
rect 19978 38904 19984 38916
rect 20036 38904 20042 38956
rect 20162 38944 20168 38956
rect 20123 38916 20168 38944
rect 20162 38904 20168 38916
rect 20220 38904 20226 38956
rect 20806 38944 20812 38956
rect 20767 38916 20812 38944
rect 20806 38904 20812 38916
rect 20864 38904 20870 38956
rect 21726 38904 21732 38956
rect 21784 38944 21790 38956
rect 22005 38947 22063 38953
rect 22005 38944 22017 38947
rect 21784 38916 22017 38944
rect 21784 38904 21790 38916
rect 22005 38913 22017 38916
rect 22051 38913 22063 38947
rect 22005 38907 22063 38913
rect 24670 38904 24676 38956
rect 24728 38944 24734 38956
rect 24780 38953 24808 38984
rect 25869 38981 25881 38984
rect 25915 38981 25927 39015
rect 31754 39012 31760 39024
rect 25869 38975 25927 38981
rect 30208 38984 31760 39012
rect 24765 38947 24823 38953
rect 24765 38944 24777 38947
rect 24728 38916 24777 38944
rect 24728 38904 24734 38916
rect 24765 38913 24777 38916
rect 24811 38913 24823 38947
rect 25038 38944 25044 38956
rect 24999 38916 25044 38944
rect 24765 38907 24823 38913
rect 25038 38904 25044 38916
rect 25096 38904 25102 38956
rect 25133 38947 25191 38953
rect 25133 38913 25145 38947
rect 25179 38913 25191 38947
rect 25133 38907 25191 38913
rect 25317 38947 25375 38953
rect 25317 38913 25329 38947
rect 25363 38944 25375 38947
rect 25406 38944 25412 38956
rect 25363 38916 25412 38944
rect 25363 38913 25375 38916
rect 25317 38907 25375 38913
rect 1854 38876 1860 38888
rect 1815 38848 1860 38876
rect 1854 38836 1860 38848
rect 1912 38836 1918 38888
rect 2041 38879 2099 38885
rect 2041 38845 2053 38879
rect 2087 38876 2099 38879
rect 2774 38876 2780 38888
rect 2087 38848 2780 38876
rect 2087 38845 2099 38848
rect 2041 38839 2099 38845
rect 2774 38836 2780 38848
rect 2832 38836 2838 38888
rect 2866 38836 2872 38888
rect 2924 38876 2930 38888
rect 14461 38879 14519 38885
rect 2924 38848 2969 38876
rect 2924 38836 2930 38848
rect 14461 38845 14473 38879
rect 14507 38876 14519 38879
rect 17037 38879 17095 38885
rect 14507 38848 16574 38876
rect 14507 38845 14519 38848
rect 14461 38839 14519 38845
rect 16546 38808 16574 38848
rect 17037 38845 17049 38879
rect 17083 38876 17095 38879
rect 17862 38876 17868 38888
rect 17083 38848 17868 38876
rect 17083 38845 17095 38848
rect 17037 38839 17095 38845
rect 17862 38836 17868 38848
rect 17920 38836 17926 38888
rect 21818 38876 21824 38888
rect 21731 38848 21824 38876
rect 21818 38836 21824 38848
rect 21876 38836 21882 38888
rect 24949 38879 25007 38885
rect 24949 38845 24961 38879
rect 24995 38845 25007 38879
rect 25148 38876 25176 38907
rect 25406 38904 25412 38916
rect 25464 38904 25470 38956
rect 25774 38944 25780 38956
rect 25735 38916 25780 38944
rect 25774 38904 25780 38916
rect 25832 38904 25838 38956
rect 26050 38944 26056 38956
rect 26011 38916 26056 38944
rect 26050 38904 26056 38916
rect 26108 38904 26114 38956
rect 30208 38953 30236 38984
rect 31754 38972 31760 38984
rect 31812 39012 31818 39024
rect 35618 39021 35624 39024
rect 35612 39012 35624 39021
rect 31812 38984 34008 39012
rect 35579 38984 35624 39012
rect 31812 38972 31818 38984
rect 33980 38956 34008 38984
rect 35612 38975 35624 38984
rect 35618 38972 35624 38975
rect 35676 38972 35682 39024
rect 30193 38947 30251 38953
rect 30193 38913 30205 38947
rect 30239 38913 30251 38947
rect 30193 38907 30251 38913
rect 30460 38947 30518 38953
rect 30460 38913 30472 38947
rect 30506 38944 30518 38947
rect 31386 38944 31392 38956
rect 30506 38916 31392 38944
rect 30506 38913 30518 38916
rect 30460 38907 30518 38913
rect 31386 38904 31392 38916
rect 31444 38904 31450 38956
rect 31846 38904 31852 38956
rect 31904 38944 31910 38956
rect 32306 38944 32312 38956
rect 31904 38916 32312 38944
rect 31904 38904 31910 38916
rect 32306 38904 32312 38916
rect 32364 38904 32370 38956
rect 33962 38904 33968 38956
rect 34020 38944 34026 38956
rect 35345 38947 35403 38953
rect 35345 38944 35357 38947
rect 34020 38916 35357 38944
rect 34020 38904 34026 38916
rect 35345 38913 35357 38916
rect 35391 38913 35403 38947
rect 37458 38944 37464 38956
rect 37419 38916 37464 38944
rect 35345 38907 35403 38913
rect 37458 38904 37464 38916
rect 37516 38904 37522 38956
rect 25222 38876 25228 38888
rect 25135 38848 25228 38876
rect 24949 38839 25007 38845
rect 21836 38808 21864 38836
rect 16546 38780 21864 38808
rect 24964 38808 24992 38839
rect 25222 38836 25228 38848
rect 25280 38876 25286 38888
rect 25792 38876 25820 38904
rect 32122 38876 32128 38888
rect 25280 38848 25820 38876
rect 32083 38848 32128 38876
rect 25280 38836 25286 38848
rect 32122 38836 32128 38848
rect 32180 38836 32186 38888
rect 25130 38808 25136 38820
rect 24964 38780 25136 38808
rect 25130 38768 25136 38780
rect 25188 38768 25194 38820
rect 34974 38768 34980 38820
rect 35032 38768 35038 38820
rect 14090 38740 14096 38752
rect 14051 38712 14096 38740
rect 14090 38700 14096 38712
rect 14148 38700 14154 38752
rect 16574 38700 16580 38752
rect 16632 38740 16638 38752
rect 16669 38743 16727 38749
rect 16669 38740 16681 38743
rect 16632 38712 16681 38740
rect 16632 38700 16638 38712
rect 16669 38709 16681 38712
rect 16715 38709 16727 38743
rect 16669 38703 16727 38709
rect 20349 38743 20407 38749
rect 20349 38709 20361 38743
rect 20395 38740 20407 38743
rect 20898 38740 20904 38752
rect 20395 38712 20904 38740
rect 20395 38709 20407 38712
rect 20349 38703 20407 38709
rect 20898 38700 20904 38712
rect 20956 38700 20962 38752
rect 23934 38700 23940 38752
rect 23992 38740 23998 38752
rect 24581 38743 24639 38749
rect 24581 38740 24593 38743
rect 23992 38712 24593 38740
rect 23992 38700 23998 38712
rect 24581 38709 24593 38712
rect 24627 38709 24639 38743
rect 24581 38703 24639 38709
rect 25866 38700 25872 38752
rect 25924 38740 25930 38752
rect 26237 38743 26295 38749
rect 26237 38740 26249 38743
rect 25924 38712 26249 38740
rect 25924 38700 25930 38712
rect 26237 38709 26249 38712
rect 26283 38709 26295 38743
rect 26237 38703 26295 38709
rect 31573 38743 31631 38749
rect 31573 38709 31585 38743
rect 31619 38740 31631 38743
rect 32306 38740 32312 38752
rect 31619 38712 32312 38740
rect 31619 38709 31631 38712
rect 31573 38703 31631 38709
rect 32306 38700 32312 38712
rect 32364 38700 32370 38752
rect 34992 38740 35020 38768
rect 36725 38743 36783 38749
rect 36725 38740 36737 38743
rect 34992 38712 36737 38740
rect 36725 38709 36737 38712
rect 36771 38709 36783 38743
rect 36725 38703 36783 38709
rect 1104 38650 38824 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 38824 38650
rect 1104 38576 38824 38598
rect 1854 38536 1860 38548
rect 1815 38508 1860 38536
rect 1854 38496 1860 38508
rect 1912 38496 1918 38548
rect 2774 38536 2780 38548
rect 2735 38508 2780 38536
rect 2774 38496 2780 38508
rect 2832 38496 2838 38548
rect 17586 38536 17592 38548
rect 17547 38508 17592 38536
rect 17586 38496 17592 38508
rect 17644 38496 17650 38548
rect 19889 38539 19947 38545
rect 19889 38505 19901 38539
rect 19935 38536 19947 38539
rect 19978 38536 19984 38548
rect 19935 38508 19984 38536
rect 19935 38505 19947 38508
rect 19889 38499 19947 38505
rect 19978 38496 19984 38508
rect 20036 38496 20042 38548
rect 20346 38536 20352 38548
rect 20307 38508 20352 38536
rect 20346 38496 20352 38508
rect 20404 38496 20410 38548
rect 32306 38536 32312 38548
rect 32267 38508 32312 38536
rect 32306 38496 32312 38508
rect 32364 38496 32370 38548
rect 18049 38471 18107 38477
rect 18049 38437 18061 38471
rect 18095 38468 18107 38471
rect 20162 38468 20168 38480
rect 18095 38440 20168 38468
rect 18095 38437 18107 38440
rect 18049 38431 18107 38437
rect 20162 38428 20168 38440
rect 20220 38428 20226 38480
rect 24854 38428 24860 38480
rect 24912 38468 24918 38480
rect 26050 38468 26056 38480
rect 24912 38440 26056 38468
rect 24912 38428 24918 38440
rect 26050 38428 26056 38440
rect 26108 38428 26114 38480
rect 17773 38403 17831 38409
rect 17773 38369 17785 38403
rect 17819 38400 17831 38403
rect 18138 38400 18144 38412
rect 17819 38372 18144 38400
rect 17819 38369 17831 38372
rect 17773 38363 17831 38369
rect 18138 38360 18144 38372
rect 18196 38400 18202 38412
rect 18598 38400 18604 38412
rect 18196 38372 18604 38400
rect 18196 38360 18202 38372
rect 18598 38360 18604 38372
rect 18656 38360 18662 38412
rect 20257 38403 20315 38409
rect 20257 38369 20269 38403
rect 20303 38400 20315 38403
rect 20346 38400 20352 38412
rect 20303 38372 20352 38400
rect 20303 38369 20315 38372
rect 20257 38363 20315 38369
rect 20346 38360 20352 38372
rect 20404 38360 20410 38412
rect 20622 38360 20628 38412
rect 20680 38400 20686 38412
rect 20680 38372 21036 38400
rect 20680 38360 20686 38372
rect 2869 38335 2927 38341
rect 2869 38301 2881 38335
rect 2915 38332 2927 38335
rect 4706 38332 4712 38344
rect 2915 38304 4712 38332
rect 2915 38301 2927 38304
rect 2869 38295 2927 38301
rect 4706 38292 4712 38304
rect 4764 38292 4770 38344
rect 15473 38335 15531 38341
rect 15473 38301 15485 38335
rect 15519 38332 15531 38335
rect 16482 38332 16488 38344
rect 15519 38304 16488 38332
rect 15519 38301 15531 38304
rect 15473 38295 15531 38301
rect 16482 38292 16488 38304
rect 16540 38292 16546 38344
rect 17862 38332 17868 38344
rect 17823 38304 17868 38332
rect 17862 38292 17868 38304
rect 17920 38292 17926 38344
rect 20070 38332 20076 38344
rect 20031 38304 20076 38332
rect 20070 38292 20076 38304
rect 20128 38332 20134 38344
rect 21008 38341 21036 38372
rect 21266 38360 21272 38412
rect 21324 38400 21330 38412
rect 22281 38403 22339 38409
rect 22281 38400 22293 38403
rect 21324 38372 22293 38400
rect 21324 38360 21330 38372
rect 22281 38369 22293 38372
rect 22327 38369 22339 38403
rect 25222 38400 25228 38412
rect 22281 38363 22339 38369
rect 24596 38372 25228 38400
rect 24596 38341 24624 38372
rect 25222 38360 25228 38372
rect 25280 38360 25286 38412
rect 32122 38360 32128 38412
rect 32180 38400 32186 38412
rect 32401 38403 32459 38409
rect 32401 38400 32413 38403
rect 32180 38372 32413 38400
rect 32180 38360 32186 38372
rect 32401 38369 32413 38372
rect 32447 38369 32459 38403
rect 37090 38400 37096 38412
rect 37051 38372 37096 38400
rect 32401 38363 32459 38369
rect 37090 38360 37096 38372
rect 37148 38360 37154 38412
rect 38105 38403 38163 38409
rect 38105 38369 38117 38403
rect 38151 38400 38163 38403
rect 38194 38400 38200 38412
rect 38151 38372 38200 38400
rect 38151 38369 38163 38372
rect 38105 38363 38163 38369
rect 38194 38360 38200 38372
rect 38252 38360 38258 38412
rect 20809 38335 20867 38341
rect 20809 38332 20821 38335
rect 20128 38304 20821 38332
rect 20128 38292 20134 38304
rect 20809 38301 20821 38304
rect 20855 38301 20867 38335
rect 20809 38295 20867 38301
rect 20993 38335 21051 38341
rect 20993 38301 21005 38335
rect 21039 38301 21051 38335
rect 20993 38295 21051 38301
rect 24581 38335 24639 38341
rect 24581 38301 24593 38335
rect 24627 38301 24639 38335
rect 24581 38295 24639 38301
rect 24670 38292 24676 38344
rect 24728 38332 24734 38344
rect 24854 38332 24860 38344
rect 24728 38304 24773 38332
rect 24815 38304 24860 38332
rect 24728 38292 24734 38304
rect 24854 38292 24860 38304
rect 24912 38292 24918 38344
rect 24949 38335 25007 38341
rect 24949 38301 24961 38335
rect 24995 38301 25007 38335
rect 24949 38295 25007 38301
rect 27433 38335 27491 38341
rect 27433 38301 27445 38335
rect 27479 38332 27491 38335
rect 27982 38332 27988 38344
rect 27479 38304 27988 38332
rect 27479 38301 27491 38304
rect 27433 38295 27491 38301
rect 15740 38267 15798 38273
rect 15740 38233 15752 38267
rect 15786 38264 15798 38267
rect 15930 38264 15936 38276
rect 15786 38236 15936 38264
rect 15786 38233 15798 38236
rect 15740 38227 15798 38233
rect 15930 38224 15936 38236
rect 15988 38224 15994 38276
rect 17589 38267 17647 38273
rect 17589 38233 17601 38267
rect 17635 38233 17647 38267
rect 17589 38227 17647 38233
rect 20349 38267 20407 38273
rect 20349 38233 20361 38267
rect 20395 38264 20407 38267
rect 20438 38264 20444 38276
rect 20395 38236 20444 38264
rect 20395 38233 20407 38236
rect 20349 38227 20407 38233
rect 16853 38199 16911 38205
rect 16853 38165 16865 38199
rect 16899 38196 16911 38199
rect 17494 38196 17500 38208
rect 16899 38168 17500 38196
rect 16899 38165 16911 38168
rect 16853 38159 16911 38165
rect 17494 38156 17500 38168
rect 17552 38196 17558 38208
rect 17604 38196 17632 38227
rect 20438 38224 20444 38236
rect 20496 38224 20502 38276
rect 22548 38267 22606 38273
rect 22548 38233 22560 38267
rect 22594 38264 22606 38267
rect 23014 38264 23020 38276
rect 22594 38236 23020 38264
rect 22594 38233 22606 38236
rect 22548 38227 22606 38233
rect 23014 38224 23020 38236
rect 23072 38224 23078 38276
rect 24964 38264 24992 38295
rect 27982 38292 27988 38304
rect 28040 38292 28046 38344
rect 30650 38292 30656 38344
rect 30708 38332 30714 38344
rect 31662 38332 31668 38344
rect 30708 38304 31668 38332
rect 30708 38292 30714 38304
rect 31662 38292 31668 38304
rect 31720 38332 31726 38344
rect 32585 38335 32643 38341
rect 32585 38332 32597 38335
rect 31720 38304 32597 38332
rect 31720 38292 31726 38304
rect 32585 38301 32597 38304
rect 32631 38301 32643 38335
rect 33594 38332 33600 38344
rect 33555 38304 33600 38332
rect 32585 38295 32643 38301
rect 33594 38292 33600 38304
rect 33652 38292 33658 38344
rect 35434 38332 35440 38344
rect 35395 38304 35440 38332
rect 35434 38292 35440 38304
rect 35492 38292 35498 38344
rect 35621 38335 35679 38341
rect 35621 38301 35633 38335
rect 35667 38332 35679 38335
rect 35894 38332 35900 38344
rect 35667 38304 35900 38332
rect 35667 38301 35679 38304
rect 35621 38295 35679 38301
rect 35894 38292 35900 38304
rect 35952 38292 35958 38344
rect 27706 38273 27712 38276
rect 23676 38236 24992 38264
rect 21174 38196 21180 38208
rect 17552 38168 17632 38196
rect 21135 38168 21180 38196
rect 17552 38156 17558 38168
rect 21174 38156 21180 38168
rect 21232 38156 21238 38208
rect 23676 38205 23704 38236
rect 24872 38208 24900 38236
rect 27700 38227 27712 38273
rect 27764 38264 27770 38276
rect 27764 38236 27800 38264
rect 27706 38224 27712 38227
rect 27764 38224 27770 38236
rect 32214 38224 32220 38276
rect 32272 38264 32278 38276
rect 32309 38267 32367 38273
rect 32309 38264 32321 38267
rect 32272 38236 32321 38264
rect 32272 38224 32278 38236
rect 32309 38233 32321 38236
rect 32355 38233 32367 38267
rect 33413 38267 33471 38273
rect 33413 38264 33425 38267
rect 32309 38227 32367 38233
rect 32784 38236 33425 38264
rect 23661 38199 23719 38205
rect 23661 38165 23673 38199
rect 23707 38165 23719 38199
rect 23661 38159 23719 38165
rect 24210 38156 24216 38208
rect 24268 38196 24274 38208
rect 24397 38199 24455 38205
rect 24397 38196 24409 38199
rect 24268 38168 24409 38196
rect 24268 38156 24274 38168
rect 24397 38165 24409 38168
rect 24443 38165 24455 38199
rect 24397 38159 24455 38165
rect 24854 38156 24860 38208
rect 24912 38156 24918 38208
rect 27522 38156 27528 38208
rect 27580 38196 27586 38208
rect 32784 38205 32812 38236
rect 33413 38233 33425 38236
rect 33459 38233 33471 38267
rect 33413 38227 33471 38233
rect 37458 38224 37464 38276
rect 37516 38264 37522 38276
rect 37921 38267 37979 38273
rect 37921 38264 37933 38267
rect 37516 38236 37933 38264
rect 37516 38224 37522 38236
rect 37921 38233 37933 38236
rect 37967 38233 37979 38267
rect 37921 38227 37979 38233
rect 28813 38199 28871 38205
rect 28813 38196 28825 38199
rect 27580 38168 28825 38196
rect 27580 38156 27586 38168
rect 28813 38165 28825 38168
rect 28859 38165 28871 38199
rect 28813 38159 28871 38165
rect 32769 38199 32827 38205
rect 32769 38165 32781 38199
rect 32815 38165 32827 38199
rect 32769 38159 32827 38165
rect 33134 38156 33140 38208
rect 33192 38196 33198 38208
rect 33229 38199 33287 38205
rect 33229 38196 33241 38199
rect 33192 38168 33241 38196
rect 33192 38156 33198 38168
rect 33229 38165 33241 38168
rect 33275 38165 33287 38199
rect 35802 38196 35808 38208
rect 35763 38168 35808 38196
rect 33229 38159 33287 38165
rect 35802 38156 35808 38168
rect 35860 38156 35866 38208
rect 1104 38106 38824 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 38824 38106
rect 1104 38032 38824 38054
rect 15930 37992 15936 38004
rect 15891 37964 15936 37992
rect 15930 37952 15936 37964
rect 15988 37952 15994 38004
rect 17770 37952 17776 38004
rect 17828 37992 17834 38004
rect 18049 37995 18107 38001
rect 18049 37992 18061 37995
rect 17828 37964 18061 37992
rect 17828 37952 17834 37964
rect 18049 37961 18061 37964
rect 18095 37992 18107 37995
rect 18138 37992 18144 38004
rect 18095 37964 18144 37992
rect 18095 37961 18107 37964
rect 18049 37955 18107 37961
rect 18138 37952 18144 37964
rect 18196 37952 18202 38004
rect 20254 37992 20260 38004
rect 20215 37964 20260 37992
rect 20254 37952 20260 37964
rect 20312 37952 20318 38004
rect 27617 37995 27675 38001
rect 27617 37961 27629 37995
rect 27663 37992 27675 37995
rect 27706 37992 27712 38004
rect 27663 37964 27712 37992
rect 27663 37961 27675 37964
rect 27617 37955 27675 37961
rect 27706 37952 27712 37964
rect 27764 37952 27770 38004
rect 29273 37995 29331 38001
rect 29273 37961 29285 37995
rect 29319 37961 29331 37995
rect 29822 37992 29828 38004
rect 29783 37964 29828 37992
rect 29273 37955 29331 37961
rect 17494 37884 17500 37936
rect 17552 37924 17558 37936
rect 20438 37924 20444 37936
rect 17552 37896 18828 37924
rect 20399 37896 20444 37924
rect 17552 37884 17558 37896
rect 14090 37856 14096 37868
rect 14051 37828 14096 37856
rect 14090 37816 14096 37828
rect 14148 37816 14154 37868
rect 16117 37859 16175 37865
rect 16117 37825 16129 37859
rect 16163 37856 16175 37859
rect 16574 37856 16580 37868
rect 16163 37828 16580 37856
rect 16163 37825 16175 37828
rect 16117 37819 16175 37825
rect 16574 37816 16580 37828
rect 16632 37816 16638 37868
rect 16758 37816 16764 37868
rect 16816 37856 16822 37868
rect 16925 37859 16983 37865
rect 16925 37856 16937 37859
rect 16816 37828 16937 37856
rect 16816 37816 16822 37828
rect 16925 37825 16937 37828
rect 16971 37825 16983 37859
rect 18690 37856 18696 37868
rect 18651 37828 18696 37856
rect 16925 37819 16983 37825
rect 18690 37816 18696 37828
rect 18748 37816 18754 37868
rect 18800 37865 18828 37896
rect 20438 37884 20444 37896
rect 20496 37884 20502 37936
rect 24854 37924 24860 37936
rect 24815 37896 24860 37924
rect 24854 37884 24860 37896
rect 24912 37884 24918 37936
rect 25314 37884 25320 37936
rect 25372 37924 25378 37936
rect 26053 37927 26111 37933
rect 26053 37924 26065 37927
rect 25372 37896 26065 37924
rect 25372 37884 25378 37896
rect 26053 37893 26065 37896
rect 26099 37893 26111 37927
rect 26053 37887 26111 37893
rect 26237 37927 26295 37933
rect 26237 37893 26249 37927
rect 26283 37924 26295 37927
rect 27522 37924 27528 37936
rect 26283 37896 27528 37924
rect 26283 37893 26295 37896
rect 26237 37887 26295 37893
rect 27522 37884 27528 37896
rect 27580 37884 27586 37936
rect 18785 37859 18843 37865
rect 18785 37825 18797 37859
rect 18831 37825 18843 37859
rect 19518 37856 19524 37868
rect 19479 37828 19524 37856
rect 18785 37819 18843 37825
rect 19518 37816 19524 37828
rect 19576 37816 19582 37868
rect 20070 37856 20076 37868
rect 20031 37828 20076 37856
rect 20070 37816 20076 37828
rect 20128 37816 20134 37868
rect 20346 37816 20352 37868
rect 20404 37856 20410 37868
rect 21085 37859 21143 37865
rect 20404 37828 20449 37856
rect 20404 37816 20410 37828
rect 21085 37825 21097 37859
rect 21131 37856 21143 37859
rect 21174 37856 21180 37868
rect 21131 37828 21180 37856
rect 21131 37825 21143 37828
rect 21085 37819 21143 37825
rect 21174 37816 21180 37828
rect 21232 37816 21238 37868
rect 23106 37856 23112 37868
rect 23067 37828 23112 37856
rect 23106 37816 23112 37828
rect 23164 37816 23170 37868
rect 23293 37859 23351 37865
rect 23293 37825 23305 37859
rect 23339 37856 23351 37859
rect 23934 37856 23940 37868
rect 23339 37828 23940 37856
rect 23339 37825 23351 37828
rect 23293 37819 23351 37825
rect 23934 37816 23940 37828
rect 23992 37816 23998 37868
rect 24118 37856 24124 37868
rect 24079 37828 24124 37856
rect 24118 37816 24124 37828
rect 24176 37816 24182 37868
rect 24210 37816 24216 37868
rect 24268 37856 24274 37868
rect 24268 37828 24313 37856
rect 24268 37816 24274 37828
rect 26786 37816 26792 37868
rect 26844 37856 26850 37868
rect 26973 37859 27031 37865
rect 26973 37856 26985 37859
rect 26844 37828 26985 37856
rect 26844 37816 26850 37828
rect 26973 37825 26985 37828
rect 27019 37825 27031 37859
rect 27157 37859 27215 37865
rect 27157 37856 27169 37859
rect 26973 37819 27031 37825
rect 27080 37828 27169 37856
rect 16482 37748 16488 37800
rect 16540 37788 16546 37800
rect 16669 37791 16727 37797
rect 16669 37788 16681 37791
rect 16540 37760 16681 37788
rect 16540 37748 16546 37760
rect 16669 37757 16681 37760
rect 16715 37757 16727 37791
rect 16669 37751 16727 37757
rect 26421 37791 26479 37797
rect 26421 37757 26433 37791
rect 26467 37788 26479 37791
rect 27080 37788 27108 37828
rect 27157 37825 27169 37828
rect 27203 37825 27215 37859
rect 27157 37819 27215 37825
rect 27249 37859 27307 37865
rect 27249 37825 27261 37859
rect 27295 37825 27307 37859
rect 27249 37819 27307 37825
rect 26467 37760 27108 37788
rect 26467 37757 26479 37760
rect 26421 37751 26479 37757
rect 27264 37732 27292 37819
rect 27338 37816 27344 37868
rect 27396 37856 27402 37868
rect 28902 37856 28908 37868
rect 27396 37828 27441 37856
rect 28863 37828 28908 37856
rect 27396 37816 27402 37828
rect 28902 37816 28908 37828
rect 28960 37816 28966 37868
rect 29288 37856 29316 37955
rect 29822 37952 29828 37964
rect 29880 37952 29886 38004
rect 32306 37952 32312 38004
rect 32364 37992 32370 38004
rect 32493 37995 32551 38001
rect 32493 37992 32505 37995
rect 32364 37964 32505 37992
rect 32364 37952 32370 37964
rect 32493 37961 32505 37964
rect 32539 37961 32551 37995
rect 37458 37992 37464 38004
rect 37419 37964 37464 37992
rect 32493 37955 32551 37961
rect 37458 37952 37464 37964
rect 37516 37952 37522 38004
rect 32122 37884 32128 37936
rect 32180 37924 32186 37936
rect 32585 37927 32643 37933
rect 32585 37924 32597 37927
rect 32180 37896 32597 37924
rect 32180 37884 32186 37896
rect 32585 37893 32597 37896
rect 32631 37893 32643 37927
rect 32585 37887 32643 37893
rect 29733 37859 29791 37865
rect 29733 37856 29745 37859
rect 29288 37828 29745 37856
rect 29733 37825 29745 37828
rect 29779 37825 29791 37859
rect 29733 37819 29791 37825
rect 30009 37859 30067 37865
rect 30009 37825 30021 37859
rect 30055 37856 30067 37859
rect 30098 37856 30104 37868
rect 30055 37828 30104 37856
rect 30055 37825 30067 37828
rect 30009 37819 30067 37825
rect 30098 37816 30104 37828
rect 30156 37816 30162 37868
rect 32214 37816 32220 37868
rect 32272 37856 32278 37868
rect 32677 37859 32735 37865
rect 32677 37856 32689 37859
rect 32272 37828 32689 37856
rect 32272 37816 32278 37828
rect 32677 37825 32689 37828
rect 32723 37825 32735 37859
rect 34514 37856 34520 37868
rect 34475 37828 34520 37856
rect 32677 37819 32735 37825
rect 34514 37816 34520 37828
rect 34572 37816 34578 37868
rect 35618 37865 35624 37868
rect 35612 37819 35624 37865
rect 35676 37856 35682 37868
rect 35676 37828 35712 37856
rect 35618 37816 35624 37819
rect 35676 37816 35682 37828
rect 37274 37816 37280 37868
rect 37332 37856 37338 37868
rect 37369 37859 37427 37865
rect 37369 37856 37381 37859
rect 37332 37828 37381 37856
rect 37332 37816 37338 37828
rect 37369 37825 37381 37828
rect 37415 37856 37427 37859
rect 38286 37856 38292 37868
rect 37415 37828 38292 37856
rect 37415 37825 37427 37828
rect 37369 37819 37427 37825
rect 38286 37816 38292 37828
rect 38344 37816 38350 37868
rect 28994 37788 29000 37800
rect 28955 37760 29000 37788
rect 28994 37748 29000 37760
rect 29052 37748 29058 37800
rect 31662 37748 31668 37800
rect 31720 37788 31726 37800
rect 32309 37791 32367 37797
rect 32309 37788 32321 37791
rect 31720 37760 32321 37788
rect 31720 37748 31726 37760
rect 32309 37757 32321 37760
rect 32355 37757 32367 37791
rect 35342 37788 35348 37800
rect 35303 37760 35348 37788
rect 32309 37751 32367 37757
rect 35342 37748 35348 37760
rect 35400 37748 35406 37800
rect 27246 37680 27252 37732
rect 27304 37680 27310 37732
rect 14277 37655 14335 37661
rect 14277 37621 14289 37655
rect 14323 37652 14335 37655
rect 14642 37652 14648 37664
rect 14323 37624 14648 37652
rect 14323 37621 14335 37624
rect 14277 37615 14335 37621
rect 14642 37612 14648 37624
rect 14700 37612 14706 37664
rect 18506 37652 18512 37664
rect 18467 37624 18512 37652
rect 18506 37612 18512 37624
rect 18564 37612 18570 37664
rect 19334 37652 19340 37664
rect 19295 37624 19340 37652
rect 19334 37612 19340 37624
rect 19392 37612 19398 37664
rect 20625 37655 20683 37661
rect 20625 37621 20637 37655
rect 20671 37652 20683 37655
rect 20714 37652 20720 37664
rect 20671 37624 20720 37652
rect 20671 37621 20683 37624
rect 20625 37615 20683 37621
rect 20714 37612 20720 37624
rect 20772 37612 20778 37664
rect 21266 37652 21272 37664
rect 21227 37624 21272 37652
rect 21266 37612 21272 37624
rect 21324 37612 21330 37664
rect 23293 37655 23351 37661
rect 23293 37621 23305 37655
rect 23339 37652 23351 37655
rect 23566 37652 23572 37664
rect 23339 37624 23572 37652
rect 23339 37621 23351 37624
rect 23293 37615 23351 37621
rect 23566 37612 23572 37624
rect 23624 37612 23630 37664
rect 23658 37612 23664 37664
rect 23716 37652 23722 37664
rect 23753 37655 23811 37661
rect 23753 37652 23765 37655
rect 23716 37624 23765 37652
rect 23716 37612 23722 37624
rect 23753 37621 23765 37624
rect 23799 37621 23811 37655
rect 24762 37652 24768 37664
rect 24723 37624 24768 37652
rect 23753 37615 23811 37621
rect 24762 37612 24768 37624
rect 24820 37652 24826 37664
rect 25406 37652 25412 37664
rect 24820 37624 25412 37652
rect 24820 37612 24826 37624
rect 25406 37612 25412 37624
rect 25464 37612 25470 37664
rect 30006 37652 30012 37664
rect 29967 37624 30012 37652
rect 30006 37612 30012 37624
rect 30064 37612 30070 37664
rect 32766 37612 32772 37664
rect 32824 37652 32830 37664
rect 32861 37655 32919 37661
rect 32861 37652 32873 37655
rect 32824 37624 32873 37652
rect 32824 37612 32830 37624
rect 32861 37621 32873 37624
rect 32907 37621 32919 37655
rect 34330 37652 34336 37664
rect 34291 37624 34336 37652
rect 32861 37615 32919 37621
rect 34330 37612 34336 37624
rect 34388 37612 34394 37664
rect 36722 37652 36728 37664
rect 36683 37624 36728 37652
rect 36722 37612 36728 37624
rect 36780 37612 36786 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 16758 37448 16764 37460
rect 16719 37420 16764 37448
rect 16758 37408 16764 37420
rect 16816 37408 16822 37460
rect 23014 37448 23020 37460
rect 22975 37420 23020 37448
rect 23014 37408 23020 37420
rect 23072 37408 23078 37460
rect 23106 37408 23112 37460
rect 23164 37448 23170 37460
rect 24581 37451 24639 37457
rect 24581 37448 24593 37451
rect 23164 37420 24593 37448
rect 23164 37408 23170 37420
rect 24581 37417 24593 37420
rect 24627 37417 24639 37451
rect 27246 37448 27252 37460
rect 27207 37420 27252 37448
rect 24581 37411 24639 37417
rect 27246 37408 27252 37420
rect 27304 37408 27310 37460
rect 28994 37448 29000 37460
rect 28955 37420 29000 37448
rect 28994 37408 29000 37420
rect 29052 37408 29058 37460
rect 34514 37408 34520 37460
rect 34572 37448 34578 37460
rect 34701 37451 34759 37457
rect 34701 37448 34713 37451
rect 34572 37420 34713 37448
rect 34572 37408 34578 37420
rect 34701 37417 34713 37420
rect 34747 37417 34759 37451
rect 35618 37448 35624 37460
rect 35579 37420 35624 37448
rect 34701 37411 34759 37417
rect 35618 37408 35624 37420
rect 35676 37408 35682 37460
rect 4706 37340 4712 37392
rect 4764 37380 4770 37392
rect 10962 37380 10968 37392
rect 4764 37352 10968 37380
rect 4764 37340 4770 37352
rect 10962 37340 10968 37352
rect 11020 37340 11026 37392
rect 17497 37383 17555 37389
rect 17497 37349 17509 37383
rect 17543 37380 17555 37383
rect 17862 37380 17868 37392
rect 17543 37352 17868 37380
rect 17543 37349 17555 37352
rect 17497 37343 17555 37349
rect 17862 37340 17868 37352
rect 17920 37340 17926 37392
rect 26237 37383 26295 37389
rect 26237 37349 26249 37383
rect 26283 37349 26295 37383
rect 26237 37343 26295 37349
rect 3326 37272 3332 37324
rect 3384 37312 3390 37324
rect 14274 37312 14280 37324
rect 3384 37284 14280 37312
rect 3384 37272 3390 37284
rect 14274 37272 14280 37284
rect 14332 37272 14338 37324
rect 18049 37315 18107 37321
rect 18049 37281 18061 37315
rect 18095 37312 18107 37315
rect 20622 37312 20628 37324
rect 18095 37284 20628 37312
rect 18095 37281 18107 37284
rect 18049 37275 18107 37281
rect 20622 37272 20628 37284
rect 20680 37272 20686 37324
rect 22830 37312 22836 37324
rect 22667 37284 22836 37312
rect 14369 37247 14427 37253
rect 14369 37213 14381 37247
rect 14415 37244 14427 37247
rect 16482 37244 16488 37256
rect 14415 37216 16488 37244
rect 14415 37213 14427 37216
rect 14369 37207 14427 37213
rect 16482 37204 16488 37216
rect 16540 37204 16546 37256
rect 16945 37247 17003 37253
rect 16945 37213 16957 37247
rect 16991 37244 17003 37247
rect 18506 37244 18512 37256
rect 16991 37216 18512 37244
rect 16991 37213 17003 37216
rect 16945 37207 17003 37213
rect 18506 37204 18512 37216
rect 18564 37204 18570 37256
rect 19426 37244 19432 37256
rect 19387 37216 19432 37244
rect 19426 37204 19432 37216
rect 19484 37204 19490 37256
rect 19613 37247 19671 37253
rect 19613 37213 19625 37247
rect 19659 37213 19671 37247
rect 19613 37207 19671 37213
rect 14642 37185 14648 37188
rect 14636 37176 14648 37185
rect 14603 37148 14648 37176
rect 14636 37139 14648 37148
rect 14642 37136 14648 37139
rect 14700 37136 14706 37188
rect 17586 37136 17592 37188
rect 17644 37176 17650 37188
rect 17681 37179 17739 37185
rect 17681 37176 17693 37179
rect 17644 37148 17693 37176
rect 17644 37136 17650 37148
rect 17681 37145 17693 37148
rect 17727 37145 17739 37179
rect 17681 37139 17739 37145
rect 17770 37136 17776 37188
rect 17828 37176 17834 37188
rect 19245 37179 19303 37185
rect 17828 37148 17873 37176
rect 17828 37136 17834 37148
rect 19245 37145 19257 37179
rect 19291 37176 19303 37179
rect 19518 37176 19524 37188
rect 19291 37148 19524 37176
rect 19291 37145 19303 37148
rect 19245 37139 19303 37145
rect 19518 37136 19524 37148
rect 19576 37136 19582 37188
rect 15749 37111 15807 37117
rect 15749 37077 15761 37111
rect 15795 37108 15807 37111
rect 16850 37108 16856 37120
rect 15795 37080 16856 37108
rect 15795 37077 15807 37080
rect 15749 37071 15807 37077
rect 16850 37068 16856 37080
rect 16908 37068 16914 37120
rect 17494 37068 17500 37120
rect 17552 37108 17558 37120
rect 17865 37111 17923 37117
rect 17865 37108 17877 37111
rect 17552 37080 17877 37108
rect 17552 37068 17558 37080
rect 17865 37077 17877 37080
rect 17911 37077 17923 37111
rect 19628 37108 19656 37207
rect 20254 37204 20260 37256
rect 20312 37244 20318 37256
rect 21913 37247 21971 37253
rect 21913 37244 21925 37247
rect 20312 37216 21925 37244
rect 20312 37204 20318 37216
rect 21913 37213 21925 37216
rect 21959 37213 21971 37247
rect 22370 37244 22376 37256
rect 22331 37216 22376 37244
rect 21913 37207 21971 37213
rect 22370 37204 22376 37216
rect 22428 37204 22434 37256
rect 22462 37204 22468 37256
rect 22520 37244 22526 37256
rect 22667 37253 22695 37284
rect 22830 37272 22836 37284
rect 22888 37272 22894 37324
rect 24762 37312 24768 37324
rect 23492 37284 24768 37312
rect 22557 37247 22615 37253
rect 22557 37244 22569 37247
rect 22520 37216 22569 37244
rect 22520 37204 22526 37216
rect 22557 37213 22569 37216
rect 22603 37213 22615 37247
rect 22557 37207 22615 37213
rect 22652 37247 22710 37253
rect 22652 37213 22664 37247
rect 22698 37213 22710 37247
rect 22652 37207 22710 37213
rect 22741 37247 22799 37253
rect 22741 37213 22753 37247
rect 22787 37244 22799 37247
rect 23492 37244 23520 37284
rect 22787 37216 23520 37244
rect 22787 37213 22799 37216
rect 22741 37207 22799 37213
rect 23566 37204 23572 37256
rect 23624 37244 23630 37256
rect 24412 37253 24440 37284
rect 24762 37272 24768 37284
rect 24820 37312 24826 37324
rect 25222 37312 25228 37324
rect 24820 37284 25228 37312
rect 24820 37272 24826 37284
rect 25222 37272 25228 37284
rect 25280 37272 25286 37324
rect 26252 37312 26280 37343
rect 27522 37340 27528 37392
rect 27580 37380 27586 37392
rect 27580 37352 27936 37380
rect 27580 37340 27586 37352
rect 26973 37315 27031 37321
rect 26252 37284 26924 37312
rect 23845 37247 23903 37253
rect 23845 37244 23857 37247
rect 23624 37216 23857 37244
rect 23624 37204 23630 37216
rect 23845 37213 23857 37216
rect 23891 37213 23903 37247
rect 23845 37207 23903 37213
rect 24397 37247 24455 37253
rect 24397 37213 24409 37247
rect 24443 37213 24455 37247
rect 24397 37207 24455 37213
rect 24581 37247 24639 37253
rect 24581 37213 24593 37247
rect 24627 37213 24639 37247
rect 24581 37207 24639 37213
rect 21266 37136 21272 37188
rect 21324 37176 21330 37188
rect 21646 37179 21704 37185
rect 21646 37176 21658 37179
rect 21324 37148 21658 37176
rect 21324 37136 21330 37148
rect 21646 37145 21658 37148
rect 21692 37145 21704 37179
rect 21646 37139 21704 37145
rect 23661 37179 23719 37185
rect 23661 37145 23673 37179
rect 23707 37176 23719 37179
rect 23750 37176 23756 37188
rect 23707 37148 23756 37176
rect 23707 37145 23719 37148
rect 23661 37139 23719 37145
rect 23750 37136 23756 37148
rect 23808 37176 23814 37188
rect 24118 37176 24124 37188
rect 23808 37148 24124 37176
rect 23808 37136 23814 37148
rect 24118 37136 24124 37148
rect 24176 37136 24182 37188
rect 24596 37176 24624 37207
rect 25314 37204 25320 37256
rect 25372 37244 25378 37256
rect 25409 37247 25467 37253
rect 25409 37244 25421 37247
rect 25372 37216 25421 37244
rect 25372 37204 25378 37216
rect 25409 37213 25421 37216
rect 25455 37213 25467 37247
rect 25409 37207 25467 37213
rect 26053 37247 26111 37253
rect 26053 37213 26065 37247
rect 26099 37213 26111 37247
rect 26234 37244 26240 37256
rect 26195 37216 26240 37244
rect 26053 37207 26111 37213
rect 25682 37176 25688 37188
rect 24596 37148 25688 37176
rect 25682 37136 25688 37148
rect 25740 37136 25746 37188
rect 26068 37176 26096 37207
rect 26234 37204 26240 37216
rect 26292 37204 26298 37256
rect 26896 37253 26924 37284
rect 26973 37281 26985 37315
rect 27019 37312 27031 37315
rect 27062 37312 27068 37324
rect 27019 37284 27068 37312
rect 27019 37281 27031 37284
rect 26973 37275 27031 37281
rect 27062 37272 27068 37284
rect 27120 37272 27126 37324
rect 27801 37315 27859 37321
rect 27801 37312 27813 37315
rect 27264 37284 27813 37312
rect 26881 37247 26939 37253
rect 26881 37213 26893 37247
rect 26927 37244 26939 37247
rect 27154 37244 27160 37256
rect 26927 37216 27160 37244
rect 26927 37213 26939 37216
rect 26881 37207 26939 37213
rect 27154 37204 27160 37216
rect 27212 37204 27218 37256
rect 27264 37176 27292 37284
rect 27801 37281 27813 37284
rect 27847 37281 27859 37315
rect 27801 37275 27859 37281
rect 27706 37244 27712 37256
rect 27667 37216 27712 37244
rect 27706 37204 27712 37216
rect 27764 37204 27770 37256
rect 27908 37253 27936 37352
rect 28537 37315 28595 37321
rect 28537 37281 28549 37315
rect 28583 37281 28595 37315
rect 28537 37275 28595 37281
rect 32033 37315 32091 37321
rect 32033 37281 32045 37315
rect 32079 37312 32091 37315
rect 32306 37312 32312 37324
rect 32079 37284 32312 37312
rect 32079 37281 32091 37284
rect 32033 37275 32091 37281
rect 27893 37247 27951 37253
rect 27893 37213 27905 37247
rect 27939 37213 27951 37247
rect 27893 37207 27951 37213
rect 26068 37148 27292 37176
rect 27724 37176 27752 37204
rect 28552 37176 28580 37275
rect 32306 37272 32312 37284
rect 32364 37272 32370 37324
rect 33226 37312 33232 37324
rect 33187 37284 33232 37312
rect 33226 37272 33232 37284
rect 33284 37272 33290 37324
rect 35069 37315 35127 37321
rect 35069 37281 35081 37315
rect 35115 37312 35127 37315
rect 36722 37312 36728 37324
rect 35115 37284 36728 37312
rect 35115 37281 35127 37284
rect 35069 37275 35127 37281
rect 36722 37272 36728 37284
rect 36780 37272 36786 37324
rect 38102 37312 38108 37324
rect 38063 37284 38108 37312
rect 38102 37272 38108 37284
rect 38160 37272 38166 37324
rect 28629 37247 28687 37253
rect 28629 37213 28641 37247
rect 28675 37244 28687 37247
rect 29549 37247 29607 37253
rect 28675 37216 29500 37244
rect 28675 37213 28687 37216
rect 28629 37207 28687 37213
rect 27724 37148 28580 37176
rect 20438 37108 20444 37120
rect 19628 37080 20444 37108
rect 17865 37071 17923 37077
rect 20438 37068 20444 37080
rect 20496 37108 20502 37120
rect 20533 37111 20591 37117
rect 20533 37108 20545 37111
rect 20496 37080 20545 37108
rect 20496 37068 20502 37080
rect 20533 37077 20545 37080
rect 20579 37077 20591 37111
rect 23474 37108 23480 37120
rect 23435 37080 23480 37108
rect 20533 37071 20591 37077
rect 23474 37068 23480 37080
rect 23532 37068 23538 37120
rect 25314 37108 25320 37120
rect 25275 37080 25320 37108
rect 25314 37068 25320 37080
rect 25372 37068 25378 37120
rect 29472 37108 29500 37216
rect 29549 37213 29561 37247
rect 29595 37244 29607 37247
rect 31754 37244 31760 37256
rect 29595 37216 31760 37244
rect 29595 37213 29607 37216
rect 29549 37207 29607 37213
rect 31754 37204 31760 37216
rect 31812 37204 31818 37256
rect 31846 37204 31852 37256
rect 31904 37244 31910 37256
rect 32766 37244 32772 37256
rect 31904 37216 31949 37244
rect 32727 37216 32772 37244
rect 31904 37204 31910 37216
rect 32766 37204 32772 37216
rect 32824 37204 32830 37256
rect 33134 37253 33140 37256
rect 33091 37247 33140 37253
rect 33091 37213 33103 37247
rect 33137 37213 33140 37247
rect 33091 37207 33140 37213
rect 33134 37204 33140 37207
rect 33192 37204 33198 37256
rect 34514 37204 34520 37256
rect 34572 37244 34578 37256
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 34572 37216 34897 37244
rect 34572 37204 34578 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 35802 37244 35808 37256
rect 35763 37216 35808 37244
rect 34885 37207 34943 37213
rect 29816 37179 29874 37185
rect 29816 37145 29828 37179
rect 29862 37176 29874 37179
rect 30006 37176 30012 37188
rect 29862 37148 30012 37176
rect 29862 37145 29874 37148
rect 29816 37139 29874 37145
rect 30006 37136 30012 37148
rect 30064 37136 30070 37188
rect 32861 37179 32919 37185
rect 32861 37145 32873 37179
rect 32907 37145 32919 37179
rect 32861 37139 32919 37145
rect 30834 37108 30840 37120
rect 29472 37080 30840 37108
rect 30834 37068 30840 37080
rect 30892 37108 30898 37120
rect 30929 37111 30987 37117
rect 30929 37108 30941 37111
rect 30892 37080 30941 37108
rect 30892 37068 30898 37080
rect 30929 37077 30941 37080
rect 30975 37077 30987 37111
rect 30929 37071 30987 37077
rect 31386 37068 31392 37120
rect 31444 37108 31450 37120
rect 31665 37111 31723 37117
rect 31665 37108 31677 37111
rect 31444 37080 31677 37108
rect 31444 37068 31450 37080
rect 31665 37077 31677 37080
rect 31711 37077 31723 37111
rect 32582 37108 32588 37120
rect 32543 37080 32588 37108
rect 31665 37071 31723 37077
rect 32582 37068 32588 37080
rect 32640 37068 32646 37120
rect 32876 37108 32904 37139
rect 32950 37136 32956 37188
rect 33008 37176 33014 37188
rect 34900 37176 34928 37207
rect 35802 37204 35808 37216
rect 35860 37204 35866 37256
rect 36262 37244 36268 37256
rect 36223 37216 36268 37244
rect 36262 37204 36268 37216
rect 36320 37204 36326 37256
rect 35986 37176 35992 37188
rect 33008 37148 33053 37176
rect 34900 37148 35992 37176
rect 33008 37136 33014 37148
rect 35986 37136 35992 37148
rect 36044 37136 36050 37188
rect 36449 37179 36507 37185
rect 36449 37145 36461 37179
rect 36495 37176 36507 37179
rect 37458 37176 37464 37188
rect 36495 37148 37464 37176
rect 36495 37145 36507 37148
rect 36449 37139 36507 37145
rect 37458 37136 37464 37148
rect 37516 37136 37522 37188
rect 34698 37108 34704 37120
rect 32876 37080 34704 37108
rect 34698 37068 34704 37080
rect 34756 37068 34762 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 19981 36907 20039 36913
rect 19981 36873 19993 36907
rect 20027 36904 20039 36907
rect 20346 36904 20352 36916
rect 20027 36876 20352 36904
rect 20027 36873 20039 36876
rect 19981 36867 20039 36873
rect 20346 36864 20352 36876
rect 20404 36864 20410 36916
rect 22462 36864 22468 36916
rect 22520 36904 22526 36916
rect 22649 36907 22707 36913
rect 22649 36904 22661 36907
rect 22520 36876 22661 36904
rect 22520 36864 22526 36876
rect 22649 36873 22661 36876
rect 22695 36873 22707 36907
rect 22649 36867 22707 36873
rect 23017 36907 23075 36913
rect 23017 36873 23029 36907
rect 23063 36904 23075 36907
rect 23474 36904 23480 36916
rect 23063 36876 23480 36904
rect 23063 36873 23075 36876
rect 23017 36867 23075 36873
rect 23474 36864 23480 36876
rect 23532 36864 23538 36916
rect 27154 36904 27160 36916
rect 27115 36876 27160 36904
rect 27154 36864 27160 36876
rect 27212 36864 27218 36916
rect 27525 36907 27583 36913
rect 27525 36873 27537 36907
rect 27571 36904 27583 36907
rect 28902 36904 28908 36916
rect 27571 36876 28908 36904
rect 27571 36873 27583 36876
rect 27525 36867 27583 36873
rect 28902 36864 28908 36876
rect 28960 36864 28966 36916
rect 30009 36907 30067 36913
rect 30009 36873 30021 36907
rect 30055 36904 30067 36907
rect 30098 36904 30104 36916
rect 30055 36876 30104 36904
rect 30055 36873 30067 36876
rect 30009 36867 30067 36873
rect 30098 36864 30104 36876
rect 30156 36864 30162 36916
rect 32122 36904 32128 36916
rect 32083 36876 32128 36904
rect 32122 36864 32128 36876
rect 32180 36864 32186 36916
rect 32766 36864 32772 36916
rect 32824 36904 32830 36916
rect 35434 36904 35440 36916
rect 32824 36876 35440 36904
rect 32824 36864 32830 36876
rect 35434 36864 35440 36876
rect 35492 36864 35498 36916
rect 37458 36904 37464 36916
rect 37419 36876 37464 36904
rect 37458 36864 37464 36876
rect 37516 36864 37522 36916
rect 14274 36836 14280 36848
rect 14235 36808 14280 36836
rect 14274 36796 14280 36808
rect 14332 36796 14338 36848
rect 20254 36836 20260 36848
rect 18616 36808 20260 36836
rect 16482 36728 16488 36780
rect 16540 36768 16546 36780
rect 18616 36777 18644 36808
rect 20254 36796 20260 36808
rect 20312 36796 20318 36848
rect 20714 36836 20720 36848
rect 20675 36808 20720 36836
rect 20714 36796 20720 36808
rect 20772 36796 20778 36848
rect 20898 36796 20904 36848
rect 20956 36845 20962 36848
rect 20956 36839 20985 36845
rect 20973 36805 20985 36839
rect 23382 36836 23388 36848
rect 20956 36799 20985 36805
rect 22848 36808 23388 36836
rect 20956 36796 20962 36799
rect 18601 36771 18659 36777
rect 18601 36768 18613 36771
rect 16540 36740 18613 36768
rect 16540 36728 16546 36740
rect 18601 36737 18613 36740
rect 18647 36737 18659 36771
rect 18601 36731 18659 36737
rect 18868 36771 18926 36777
rect 18868 36737 18880 36771
rect 18914 36768 18926 36771
rect 19334 36768 19340 36780
rect 18914 36740 19340 36768
rect 18914 36737 18926 36740
rect 18868 36731 18926 36737
rect 19334 36728 19340 36740
rect 19392 36728 19398 36780
rect 20622 36768 20628 36780
rect 20583 36740 20628 36768
rect 20622 36728 20628 36740
rect 20680 36728 20686 36780
rect 22848 36777 22876 36808
rect 23382 36796 23388 36808
rect 23440 36796 23446 36848
rect 25406 36796 25412 36848
rect 25464 36836 25470 36848
rect 26053 36839 26111 36845
rect 26053 36836 26065 36839
rect 25464 36808 26065 36836
rect 25464 36796 25470 36808
rect 26053 36805 26065 36808
rect 26099 36805 26111 36839
rect 26053 36799 26111 36805
rect 26234 36796 26240 36848
rect 26292 36836 26298 36848
rect 26970 36836 26976 36848
rect 26292 36808 26976 36836
rect 26292 36796 26298 36808
rect 26970 36796 26976 36808
rect 27028 36836 27034 36848
rect 27028 36808 27384 36836
rect 27028 36796 27034 36808
rect 20809 36771 20867 36777
rect 20809 36737 20821 36771
rect 20855 36737 20867 36771
rect 20809 36731 20867 36737
rect 22833 36771 22891 36777
rect 22833 36737 22845 36771
rect 22879 36737 22891 36771
rect 22833 36731 22891 36737
rect 23109 36771 23167 36777
rect 23109 36737 23121 36771
rect 23155 36737 23167 36771
rect 23566 36768 23572 36780
rect 23527 36740 23572 36768
rect 23109 36731 23167 36737
rect 14366 36660 14372 36712
rect 14424 36700 14430 36712
rect 15933 36703 15991 36709
rect 15933 36700 15945 36703
rect 14424 36672 15945 36700
rect 14424 36660 14430 36672
rect 15933 36669 15945 36672
rect 15979 36669 15991 36703
rect 15933 36663 15991 36669
rect 16117 36703 16175 36709
rect 16117 36669 16129 36703
rect 16163 36669 16175 36703
rect 16117 36663 16175 36669
rect 15746 36592 15752 36644
rect 15804 36632 15810 36644
rect 16132 36632 16160 36663
rect 20714 36660 20720 36712
rect 20772 36700 20778 36712
rect 20824 36700 20852 36731
rect 21085 36703 21143 36709
rect 21085 36700 21097 36703
rect 20772 36672 20852 36700
rect 20916 36672 21097 36700
rect 20772 36660 20778 36672
rect 20916 36644 20944 36672
rect 21085 36669 21097 36672
rect 21131 36669 21143 36703
rect 23124 36700 23152 36731
rect 23566 36728 23572 36740
rect 23624 36728 23630 36780
rect 23750 36768 23756 36780
rect 23711 36740 23756 36768
rect 23750 36728 23756 36740
rect 23808 36728 23814 36780
rect 24946 36728 24952 36780
rect 25004 36768 25010 36780
rect 25314 36768 25320 36780
rect 25004 36740 25320 36768
rect 25004 36728 25010 36740
rect 25314 36728 25320 36740
rect 25372 36728 25378 36780
rect 27062 36768 27068 36780
rect 27023 36740 27068 36768
rect 27062 36728 27068 36740
rect 27120 36728 27126 36780
rect 27356 36777 27384 36808
rect 30742 36796 30748 36848
rect 30800 36836 30806 36848
rect 31113 36839 31171 36845
rect 31113 36836 31125 36839
rect 30800 36808 31125 36836
rect 30800 36796 30806 36808
rect 31113 36805 31125 36808
rect 31159 36805 31171 36839
rect 31113 36799 31171 36805
rect 31297 36839 31355 36845
rect 31297 36805 31309 36839
rect 31343 36836 31355 36839
rect 31754 36836 31760 36848
rect 31343 36808 31760 36836
rect 31343 36805 31355 36808
rect 31297 36799 31355 36805
rect 31754 36796 31760 36808
rect 31812 36836 31818 36848
rect 32858 36836 32864 36848
rect 31812 36808 32864 36836
rect 31812 36796 31818 36808
rect 32858 36796 32864 36808
rect 32916 36796 32922 36848
rect 34232 36839 34290 36845
rect 34232 36805 34244 36839
rect 34278 36836 34290 36839
rect 34330 36836 34336 36848
rect 34278 36808 34336 36836
rect 34278 36805 34290 36808
rect 34232 36799 34290 36805
rect 34330 36796 34336 36808
rect 34388 36796 34394 36848
rect 27341 36771 27399 36777
rect 27341 36737 27353 36771
rect 27387 36737 27399 36771
rect 27341 36731 27399 36737
rect 29733 36771 29791 36777
rect 29733 36737 29745 36771
rect 29779 36768 29791 36771
rect 30834 36768 30840 36780
rect 29779 36740 30840 36768
rect 29779 36737 29791 36740
rect 29733 36731 29791 36737
rect 30834 36728 30840 36740
rect 30892 36728 30898 36780
rect 31570 36728 31576 36780
rect 31628 36768 31634 36780
rect 33238 36771 33296 36777
rect 33238 36768 33250 36771
rect 31628 36740 33250 36768
rect 31628 36728 31634 36740
rect 33238 36737 33250 36740
rect 33284 36737 33296 36771
rect 33238 36731 33296 36737
rect 36262 36728 36268 36780
rect 36320 36768 36326 36780
rect 36541 36771 36599 36777
rect 36541 36768 36553 36771
rect 36320 36740 36553 36768
rect 36320 36728 36326 36740
rect 36541 36737 36553 36740
rect 36587 36737 36599 36771
rect 37366 36768 37372 36780
rect 37279 36740 37372 36768
rect 36541 36731 36599 36737
rect 37366 36728 37372 36740
rect 37424 36768 37430 36780
rect 38470 36768 38476 36780
rect 37424 36740 38476 36768
rect 37424 36728 37430 36740
rect 38470 36728 38476 36740
rect 38528 36728 38534 36780
rect 23661 36703 23719 36709
rect 23661 36700 23673 36703
rect 23124 36672 23673 36700
rect 21085 36663 21143 36669
rect 23661 36669 23673 36672
rect 23707 36669 23719 36703
rect 23661 36663 23719 36669
rect 29546 36660 29552 36712
rect 29604 36700 29610 36712
rect 30009 36703 30067 36709
rect 30009 36700 30021 36703
rect 29604 36672 30021 36700
rect 29604 36660 29610 36672
rect 30009 36669 30021 36672
rect 30055 36700 30067 36703
rect 30190 36700 30196 36712
rect 30055 36672 30196 36700
rect 30055 36669 30067 36672
rect 30009 36663 30067 36669
rect 30190 36660 30196 36672
rect 30248 36660 30254 36712
rect 33505 36703 33563 36709
rect 33505 36669 33517 36703
rect 33551 36700 33563 36703
rect 33965 36703 34023 36709
rect 33965 36700 33977 36703
rect 33551 36672 33977 36700
rect 33551 36669 33563 36672
rect 33505 36663 33563 36669
rect 33965 36669 33977 36672
rect 34011 36669 34023 36703
rect 33965 36663 34023 36669
rect 15804 36604 16160 36632
rect 15804 36592 15810 36604
rect 20898 36592 20904 36644
rect 20956 36592 20962 36644
rect 26050 36592 26056 36644
rect 26108 36632 26114 36644
rect 26237 36635 26295 36641
rect 26237 36632 26249 36635
rect 26108 36604 26249 36632
rect 26108 36592 26114 36604
rect 26237 36601 26249 36604
rect 26283 36632 26295 36635
rect 29638 36632 29644 36644
rect 26283 36604 29644 36632
rect 26283 36601 26295 36604
rect 26237 36595 26295 36601
rect 29638 36592 29644 36604
rect 29696 36632 29702 36644
rect 29825 36635 29883 36641
rect 29825 36632 29837 36635
rect 29696 36604 29837 36632
rect 29696 36592 29702 36604
rect 29825 36601 29837 36604
rect 29871 36601 29883 36635
rect 29825 36595 29883 36601
rect 20438 36564 20444 36576
rect 20399 36536 20444 36564
rect 20438 36524 20444 36536
rect 20496 36524 20502 36576
rect 23382 36524 23388 36576
rect 23440 36564 23446 36576
rect 25409 36567 25467 36573
rect 25409 36564 25421 36567
rect 23440 36536 25421 36564
rect 23440 36524 23446 36536
rect 25409 36533 25421 36536
rect 25455 36564 25467 36567
rect 26602 36564 26608 36576
rect 25455 36536 26608 36564
rect 25455 36533 25467 36536
rect 25409 36527 25467 36533
rect 26602 36524 26608 36536
rect 26660 36564 26666 36576
rect 27338 36564 27344 36576
rect 26660 36536 27344 36564
rect 26660 36524 26666 36536
rect 27338 36524 27344 36536
rect 27396 36524 27402 36576
rect 30190 36524 30196 36576
rect 30248 36564 30254 36576
rect 32766 36564 32772 36576
rect 30248 36536 32772 36564
rect 30248 36524 30254 36536
rect 32766 36524 32772 36536
rect 32824 36524 32830 36576
rect 32858 36524 32864 36576
rect 32916 36564 32922 36576
rect 33520 36564 33548 36663
rect 32916 36536 33548 36564
rect 32916 36524 32922 36536
rect 34606 36524 34612 36576
rect 34664 36564 34670 36576
rect 35345 36567 35403 36573
rect 35345 36564 35357 36567
rect 34664 36536 35357 36564
rect 34664 36524 34670 36536
rect 35345 36533 35357 36536
rect 35391 36533 35403 36567
rect 35345 36527 35403 36533
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 14366 36360 14372 36372
rect 14327 36332 14372 36360
rect 14366 36320 14372 36332
rect 14424 36320 14430 36372
rect 20254 36360 20260 36372
rect 20215 36332 20260 36360
rect 20254 36320 20260 36332
rect 20312 36320 20318 36372
rect 37366 36360 37372 36372
rect 20364 36332 37372 36360
rect 19242 36252 19248 36304
rect 19300 36292 19306 36304
rect 20364 36292 20392 36332
rect 37366 36320 37372 36332
rect 37424 36320 37430 36372
rect 19300 36264 20392 36292
rect 19300 36252 19306 36264
rect 21634 36252 21640 36304
rect 21692 36292 21698 36304
rect 21729 36295 21787 36301
rect 21729 36292 21741 36295
rect 21692 36264 21741 36292
rect 21692 36252 21698 36264
rect 21729 36261 21741 36264
rect 21775 36292 21787 36295
rect 22370 36292 22376 36304
rect 21775 36264 22376 36292
rect 21775 36261 21787 36264
rect 21729 36255 21787 36261
rect 22370 36252 22376 36264
rect 22428 36252 22434 36304
rect 24670 36292 24676 36304
rect 24631 36264 24676 36292
rect 24670 36252 24676 36264
rect 24728 36252 24734 36304
rect 26970 36292 26976 36304
rect 26931 36264 26976 36292
rect 26970 36252 26976 36264
rect 27028 36252 27034 36304
rect 31570 36292 31576 36304
rect 31531 36264 31576 36292
rect 31570 36252 31576 36264
rect 31628 36252 31634 36304
rect 21082 36224 21088 36236
rect 20364 36196 21088 36224
rect 1394 36156 1400 36168
rect 1355 36128 1400 36156
rect 1394 36116 1400 36128
rect 1452 36116 1458 36168
rect 3234 36116 3240 36168
rect 3292 36156 3298 36168
rect 3292 36128 3337 36156
rect 3292 36116 3298 36128
rect 14090 36116 14096 36168
rect 14148 36156 14154 36168
rect 20364 36165 20392 36196
rect 21082 36184 21088 36196
rect 21140 36224 21146 36236
rect 26234 36224 26240 36236
rect 21140 36196 26240 36224
rect 21140 36184 21146 36196
rect 26234 36184 26240 36196
rect 26292 36184 26298 36236
rect 14277 36159 14335 36165
rect 14277 36156 14289 36159
rect 14148 36128 14289 36156
rect 14148 36116 14154 36128
rect 14277 36125 14289 36128
rect 14323 36125 14335 36159
rect 14277 36119 14335 36125
rect 20349 36159 20407 36165
rect 20349 36125 20361 36159
rect 20395 36125 20407 36159
rect 20349 36119 20407 36125
rect 21545 36159 21603 36165
rect 21545 36125 21557 36159
rect 21591 36156 21603 36159
rect 21818 36156 21824 36168
rect 21591 36128 21824 36156
rect 21591 36125 21603 36128
rect 21545 36119 21603 36125
rect 21818 36116 21824 36128
rect 21876 36156 21882 36168
rect 23842 36156 23848 36168
rect 21876 36128 23848 36156
rect 21876 36116 21882 36128
rect 23842 36116 23848 36128
rect 23900 36116 23906 36168
rect 24394 36156 24400 36168
rect 24355 36128 24400 36156
rect 24394 36116 24400 36128
rect 24452 36116 24458 36168
rect 25866 36156 25872 36168
rect 25827 36128 25872 36156
rect 25866 36116 25872 36128
rect 25924 36116 25930 36168
rect 26053 36159 26111 36165
rect 26053 36125 26065 36159
rect 26099 36156 26111 36159
rect 27154 36156 27160 36168
rect 26099 36128 27160 36156
rect 26099 36125 26111 36128
rect 26053 36119 26111 36125
rect 27154 36116 27160 36128
rect 27212 36116 27218 36168
rect 27341 36159 27399 36165
rect 27341 36125 27353 36159
rect 27387 36156 27399 36159
rect 27522 36156 27528 36168
rect 27387 36128 27528 36156
rect 27387 36125 27399 36128
rect 27341 36119 27399 36125
rect 27522 36116 27528 36128
rect 27580 36156 27586 36168
rect 29270 36156 29276 36168
rect 27580 36128 29276 36156
rect 27580 36116 27586 36128
rect 29270 36116 29276 36128
rect 29328 36116 29334 36168
rect 31386 36156 31392 36168
rect 31347 36128 31392 36156
rect 31386 36116 31392 36128
rect 31444 36116 31450 36168
rect 35342 36116 35348 36168
rect 35400 36156 35406 36168
rect 36170 36156 36176 36168
rect 35400 36128 36176 36156
rect 35400 36116 35406 36128
rect 36170 36116 36176 36128
rect 36228 36156 36234 36168
rect 36265 36159 36323 36165
rect 36265 36156 36277 36159
rect 36228 36128 36277 36156
rect 36228 36116 36234 36128
rect 36265 36125 36277 36128
rect 36311 36125 36323 36159
rect 36265 36119 36323 36125
rect 3050 36088 3056 36100
rect 3011 36060 3056 36088
rect 3050 36048 3056 36060
rect 3108 36048 3114 36100
rect 24578 36048 24584 36100
rect 24636 36088 24642 36100
rect 24673 36091 24731 36097
rect 24673 36088 24685 36091
rect 24636 36060 24685 36088
rect 24636 36048 24642 36060
rect 24673 36057 24685 36060
rect 24719 36057 24731 36091
rect 24673 36051 24731 36057
rect 36354 36048 36360 36100
rect 36412 36088 36418 36100
rect 36510 36091 36568 36097
rect 36510 36088 36522 36091
rect 36412 36060 36522 36088
rect 36412 36048 36418 36060
rect 36510 36057 36522 36060
rect 36556 36057 36568 36091
rect 36510 36051 36568 36057
rect 20714 35980 20720 36032
rect 20772 36020 20778 36032
rect 24302 36020 24308 36032
rect 20772 35992 24308 36020
rect 20772 35980 20778 35992
rect 24302 35980 24308 35992
rect 24360 35980 24366 36032
rect 24489 36023 24547 36029
rect 24489 35989 24501 36023
rect 24535 36020 24547 36023
rect 24854 36020 24860 36032
rect 24535 35992 24860 36020
rect 24535 35989 24547 35992
rect 24489 35983 24547 35989
rect 24854 35980 24860 35992
rect 24912 35980 24918 36032
rect 37458 35980 37464 36032
rect 37516 36020 37522 36032
rect 37645 36023 37703 36029
rect 37645 36020 37657 36023
rect 37516 35992 37657 36020
rect 37516 35980 37522 35992
rect 37645 35989 37657 35992
rect 37691 35989 37703 36023
rect 37645 35983 37703 35989
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 2777 35819 2835 35825
rect 2777 35785 2789 35819
rect 2823 35816 2835 35819
rect 3050 35816 3056 35828
rect 2823 35788 3056 35816
rect 2823 35785 2835 35788
rect 2777 35779 2835 35785
rect 3050 35776 3056 35788
rect 3108 35776 3114 35828
rect 24026 35776 24032 35828
rect 24084 35816 24090 35828
rect 36173 35819 36231 35825
rect 24084 35788 31754 35816
rect 24084 35776 24090 35788
rect 20156 35751 20214 35757
rect 20156 35717 20168 35751
rect 20202 35748 20214 35751
rect 20438 35748 20444 35760
rect 20202 35720 20444 35748
rect 20202 35717 20214 35720
rect 20156 35711 20214 35717
rect 20438 35708 20444 35720
rect 20496 35708 20502 35760
rect 23293 35751 23351 35757
rect 23293 35717 23305 35751
rect 23339 35748 23351 35751
rect 23658 35748 23664 35760
rect 23339 35720 23664 35748
rect 23339 35717 23351 35720
rect 23293 35711 23351 35717
rect 23658 35708 23664 35720
rect 23716 35708 23722 35760
rect 24486 35708 24492 35760
rect 24544 35748 24550 35760
rect 24544 35720 25544 35748
rect 24544 35708 24550 35720
rect 2869 35683 2927 35689
rect 2869 35649 2881 35683
rect 2915 35680 2927 35683
rect 14090 35680 14096 35692
rect 2915 35652 14096 35680
rect 2915 35649 2927 35652
rect 2869 35643 2927 35649
rect 14090 35640 14096 35652
rect 14148 35640 14154 35692
rect 17402 35680 17408 35692
rect 17363 35652 17408 35680
rect 17402 35640 17408 35652
rect 17460 35640 17466 35692
rect 23106 35680 23112 35692
rect 23067 35652 23112 35680
rect 23106 35640 23112 35652
rect 23164 35640 23170 35692
rect 23842 35640 23848 35692
rect 23900 35680 23906 35692
rect 24394 35680 24400 35692
rect 23900 35652 24400 35680
rect 23900 35640 23906 35652
rect 24394 35640 24400 35652
rect 24452 35680 24458 35692
rect 24765 35683 24823 35689
rect 24765 35680 24777 35683
rect 24452 35652 24777 35680
rect 24452 35640 24458 35652
rect 24765 35649 24777 35652
rect 24811 35649 24823 35683
rect 24946 35680 24952 35692
rect 24907 35652 24952 35680
rect 24765 35643 24823 35649
rect 24946 35640 24952 35652
rect 25004 35640 25010 35692
rect 25516 35689 25544 35720
rect 27154 35708 27160 35760
rect 27212 35748 27218 35760
rect 27433 35751 27491 35757
rect 27433 35748 27445 35751
rect 27212 35720 27445 35748
rect 27212 35708 27218 35720
rect 27433 35717 27445 35720
rect 27479 35748 27491 35751
rect 28074 35748 28080 35760
rect 27479 35720 28080 35748
rect 27479 35717 27491 35720
rect 27433 35711 27491 35717
rect 28074 35708 28080 35720
rect 28132 35708 28138 35760
rect 31726 35748 31754 35788
rect 36173 35785 36185 35819
rect 36219 35816 36231 35819
rect 36354 35816 36360 35828
rect 36219 35788 36360 35816
rect 36219 35785 36231 35788
rect 36173 35779 36231 35785
rect 36354 35776 36360 35788
rect 36412 35776 36418 35828
rect 31726 35720 37872 35748
rect 25501 35683 25559 35689
rect 25501 35649 25513 35683
rect 25547 35649 25559 35683
rect 25682 35680 25688 35692
rect 25643 35652 25688 35680
rect 25501 35643 25559 35649
rect 25682 35640 25688 35652
rect 25740 35680 25746 35692
rect 27617 35683 27675 35689
rect 27617 35680 27629 35683
rect 25740 35652 27629 35680
rect 25740 35640 25746 35652
rect 27617 35649 27629 35652
rect 27663 35680 27675 35683
rect 27706 35680 27712 35692
rect 27663 35652 27712 35680
rect 27663 35649 27675 35652
rect 27617 35643 27675 35649
rect 27706 35640 27712 35652
rect 27764 35640 27770 35692
rect 33413 35683 33471 35689
rect 33413 35649 33425 35683
rect 33459 35680 33471 35683
rect 33873 35683 33931 35689
rect 33873 35680 33885 35683
rect 33459 35652 33885 35680
rect 33459 35649 33471 35652
rect 33413 35643 33471 35649
rect 33873 35649 33885 35652
rect 33919 35649 33931 35683
rect 33873 35643 33931 35649
rect 34057 35683 34115 35689
rect 34057 35649 34069 35683
rect 34103 35680 34115 35683
rect 34514 35680 34520 35692
rect 34103 35652 34520 35680
rect 34103 35649 34115 35652
rect 34057 35643 34115 35649
rect 34514 35640 34520 35652
rect 34572 35640 34578 35692
rect 34698 35680 34704 35692
rect 34659 35652 34704 35680
rect 34698 35640 34704 35652
rect 34756 35640 34762 35692
rect 35989 35683 36047 35689
rect 35989 35649 36001 35683
rect 36035 35680 36047 35683
rect 36538 35680 36544 35692
rect 36035 35652 36544 35680
rect 36035 35649 36047 35652
rect 35989 35643 36047 35649
rect 36538 35640 36544 35652
rect 36596 35640 36602 35692
rect 37844 35689 37872 35720
rect 37829 35683 37887 35689
rect 37829 35649 37841 35683
rect 37875 35649 37887 35683
rect 37829 35643 37887 35649
rect 2133 35615 2191 35621
rect 2133 35581 2145 35615
rect 2179 35612 2191 35615
rect 3234 35612 3240 35624
rect 2179 35584 3240 35612
rect 2179 35581 2191 35584
rect 2133 35575 2191 35581
rect 3234 35572 3240 35584
rect 3292 35572 3298 35624
rect 19889 35615 19947 35621
rect 19889 35581 19901 35615
rect 19935 35581 19947 35615
rect 19889 35575 19947 35581
rect 17218 35476 17224 35488
rect 17179 35448 17224 35476
rect 17218 35436 17224 35448
rect 17276 35436 17282 35488
rect 19904 35476 19932 35575
rect 24578 35572 24584 35624
rect 24636 35612 24642 35624
rect 24673 35615 24731 35621
rect 24673 35612 24685 35615
rect 24636 35584 24685 35612
rect 24636 35572 24642 35584
rect 24673 35581 24685 35584
rect 24719 35581 24731 35615
rect 24673 35575 24731 35581
rect 24854 35572 24860 35624
rect 24912 35612 24918 35624
rect 25593 35615 25651 35621
rect 25593 35612 25605 35615
rect 24912 35584 25605 35612
rect 24912 35572 24918 35584
rect 25593 35581 25605 35584
rect 25639 35581 25651 35615
rect 25593 35575 25651 35581
rect 33778 35572 33784 35624
rect 33836 35612 33842 35624
rect 34241 35615 34299 35621
rect 34241 35612 34253 35615
rect 33836 35584 34253 35612
rect 33836 35572 33842 35584
rect 34241 35581 34253 35584
rect 34287 35612 34299 35615
rect 34606 35612 34612 35624
rect 34287 35584 34612 35612
rect 34287 35581 34299 35584
rect 34241 35575 34299 35581
rect 34606 35572 34612 35584
rect 34664 35612 34670 35624
rect 35434 35612 35440 35624
rect 34664 35584 35440 35612
rect 34664 35572 34670 35584
rect 35434 35572 35440 35584
rect 35492 35572 35498 35624
rect 38102 35612 38108 35624
rect 38063 35584 38108 35612
rect 38102 35572 38108 35584
rect 38160 35572 38166 35624
rect 24302 35504 24308 35556
rect 24360 35544 24366 35556
rect 30650 35544 30656 35556
rect 24360 35516 30656 35544
rect 24360 35504 24366 35516
rect 30650 35504 30656 35516
rect 30708 35504 30714 35556
rect 20162 35476 20168 35488
rect 19904 35448 20168 35476
rect 20162 35436 20168 35448
rect 20220 35436 20226 35488
rect 21266 35476 21272 35488
rect 21227 35448 21272 35476
rect 21266 35436 21272 35448
rect 21324 35436 21330 35488
rect 23477 35479 23535 35485
rect 23477 35445 23489 35479
rect 23523 35476 23535 35479
rect 23750 35476 23756 35488
rect 23523 35448 23756 35476
rect 23523 35445 23535 35448
rect 23477 35439 23535 35445
rect 23750 35436 23756 35448
rect 23808 35436 23814 35488
rect 24489 35479 24547 35485
rect 24489 35445 24501 35479
rect 24535 35476 24547 35479
rect 24762 35476 24768 35488
rect 24535 35448 24768 35476
rect 24535 35445 24547 35448
rect 24489 35439 24547 35445
rect 24762 35436 24768 35448
rect 24820 35436 24826 35488
rect 24854 35436 24860 35488
rect 24912 35476 24918 35488
rect 25866 35476 25872 35488
rect 24912 35448 25872 35476
rect 24912 35436 24918 35448
rect 25866 35436 25872 35448
rect 25924 35436 25930 35488
rect 33226 35476 33232 35488
rect 33187 35448 33232 35476
rect 33226 35436 33232 35448
rect 33284 35436 33290 35488
rect 34790 35436 34796 35488
rect 34848 35476 34854 35488
rect 34885 35479 34943 35485
rect 34885 35476 34897 35479
rect 34848 35448 34897 35476
rect 34848 35436 34854 35448
rect 34885 35445 34897 35448
rect 34931 35445 34943 35479
rect 34885 35439 34943 35445
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 17402 35272 17408 35284
rect 17363 35244 17408 35272
rect 17402 35232 17408 35244
rect 17460 35232 17466 35284
rect 20809 35275 20867 35281
rect 20809 35241 20821 35275
rect 20855 35272 20867 35275
rect 20898 35272 20904 35284
rect 20855 35244 20904 35272
rect 20855 35241 20867 35244
rect 20809 35235 20867 35241
rect 20898 35232 20904 35244
rect 20956 35232 20962 35284
rect 24854 35272 24860 35284
rect 22848 35244 24860 35272
rect 22649 35139 22707 35145
rect 17604 35108 18460 35136
rect 15562 35068 15568 35080
rect 15523 35040 15568 35068
rect 15562 35028 15568 35040
rect 15620 35028 15626 35080
rect 17604 35077 17632 35108
rect 17589 35071 17647 35077
rect 17589 35037 17601 35071
rect 17635 35037 17647 35071
rect 17589 35031 17647 35037
rect 17681 35071 17739 35077
rect 17681 35037 17693 35071
rect 17727 35037 17739 35071
rect 18322 35068 18328 35080
rect 18283 35040 18328 35068
rect 17681 35031 17739 35037
rect 15832 35003 15890 35009
rect 15832 34969 15844 35003
rect 15878 35000 15890 35003
rect 15930 35000 15936 35012
rect 15878 34972 15936 35000
rect 15878 34969 15890 34972
rect 15832 34963 15890 34969
rect 15930 34960 15936 34972
rect 15988 34960 15994 35012
rect 17696 35000 17724 35031
rect 18322 35028 18328 35040
rect 18380 35028 18386 35080
rect 18432 35077 18460 35108
rect 22649 35105 22661 35139
rect 22695 35136 22707 35139
rect 22848 35136 22876 35244
rect 24854 35232 24860 35244
rect 24912 35232 24918 35284
rect 25056 35244 26004 35272
rect 23382 35164 23388 35216
rect 23440 35204 23446 35216
rect 23440 35176 23612 35204
rect 23440 35164 23446 35176
rect 22695 35108 22876 35136
rect 22925 35139 22983 35145
rect 22695 35105 22707 35108
rect 22649 35099 22707 35105
rect 22925 35105 22937 35139
rect 22971 35105 22983 35139
rect 22925 35099 22983 35105
rect 18417 35071 18475 35077
rect 18417 35037 18429 35071
rect 18463 35068 18475 35071
rect 18690 35068 18696 35080
rect 18463 35040 18696 35068
rect 18463 35037 18475 35040
rect 18417 35031 18475 35037
rect 18690 35028 18696 35040
rect 18748 35028 18754 35080
rect 20625 35071 20683 35077
rect 20625 35037 20637 35071
rect 20671 35068 20683 35071
rect 20806 35068 20812 35080
rect 20671 35040 20812 35068
rect 20671 35037 20683 35040
rect 20625 35031 20683 35037
rect 20806 35028 20812 35040
rect 20864 35028 20870 35080
rect 22557 35071 22615 35077
rect 22557 35037 22569 35071
rect 22603 35068 22615 35071
rect 22738 35068 22744 35080
rect 22603 35040 22744 35068
rect 22603 35037 22615 35040
rect 22557 35031 22615 35037
rect 22738 35028 22744 35040
rect 22796 35028 22802 35080
rect 17862 35000 17868 35012
rect 16960 34972 17868 35000
rect 16960 34941 16988 34972
rect 17862 34960 17868 34972
rect 17920 34960 17926 35012
rect 22940 35000 22968 35099
rect 23584 35077 23612 35176
rect 23750 35164 23756 35216
rect 23808 35164 23814 35216
rect 24578 35204 24584 35216
rect 24491 35176 24584 35204
rect 24578 35164 24584 35176
rect 24636 35204 24642 35216
rect 25056 35204 25084 35244
rect 24636 35176 25084 35204
rect 24636 35164 24642 35176
rect 23768 35077 23796 35164
rect 24854 35136 24860 35148
rect 24815 35108 24860 35136
rect 24854 35096 24860 35108
rect 24912 35096 24918 35148
rect 25774 35136 25780 35148
rect 25735 35108 25780 35136
rect 25774 35096 25780 35108
rect 25832 35096 25838 35148
rect 25976 35145 26004 35244
rect 27062 35232 27068 35284
rect 27120 35272 27126 35284
rect 27709 35275 27767 35281
rect 27709 35272 27721 35275
rect 27120 35244 27721 35272
rect 27120 35232 27126 35244
rect 27709 35241 27721 35244
rect 27755 35241 27767 35275
rect 36538 35272 36544 35284
rect 36499 35244 36544 35272
rect 27709 35235 27767 35241
rect 36538 35232 36544 35244
rect 36596 35232 36602 35284
rect 26418 35164 26424 35216
rect 26476 35204 26482 35216
rect 26697 35207 26755 35213
rect 26697 35204 26709 35207
rect 26476 35176 26709 35204
rect 26476 35164 26482 35176
rect 26697 35173 26709 35176
rect 26743 35204 26755 35207
rect 36081 35207 36139 35213
rect 26743 35176 27568 35204
rect 26743 35173 26755 35176
rect 26697 35167 26755 35173
rect 25961 35139 26019 35145
rect 25961 35105 25973 35139
rect 26007 35105 26019 35139
rect 27154 35136 27160 35148
rect 27115 35108 27160 35136
rect 25961 35099 26019 35105
rect 27154 35096 27160 35108
rect 27212 35096 27218 35148
rect 27540 35080 27568 35176
rect 36081 35173 36093 35207
rect 36127 35173 36139 35207
rect 36081 35167 36139 35173
rect 27893 35139 27951 35145
rect 27893 35105 27905 35139
rect 27939 35136 27951 35139
rect 29546 35136 29552 35148
rect 27939 35108 29552 35136
rect 27939 35105 27951 35108
rect 27893 35099 27951 35105
rect 29546 35096 29552 35108
rect 29604 35096 29610 35148
rect 29638 35096 29644 35148
rect 29696 35136 29702 35148
rect 30009 35139 30067 35145
rect 30009 35136 30021 35139
rect 29696 35108 30021 35136
rect 29696 35096 29702 35108
rect 30009 35105 30021 35108
rect 30055 35105 30067 35139
rect 30190 35136 30196 35148
rect 30151 35108 30196 35136
rect 30009 35099 30067 35105
rect 30190 35096 30196 35108
rect 30248 35096 30254 35148
rect 36096 35136 36124 35167
rect 36354 35136 36360 35148
rect 36096 35108 36360 35136
rect 36354 35096 36360 35108
rect 36412 35136 36418 35148
rect 36909 35139 36967 35145
rect 36909 35136 36921 35139
rect 36412 35108 36921 35136
rect 36412 35096 36418 35108
rect 36909 35105 36921 35108
rect 36955 35105 36967 35139
rect 36909 35099 36967 35105
rect 23569 35071 23627 35077
rect 23569 35037 23581 35071
rect 23615 35037 23627 35071
rect 23569 35031 23627 35037
rect 23753 35071 23811 35077
rect 23753 35037 23765 35071
rect 23799 35037 23811 35071
rect 23753 35031 23811 35037
rect 23842 35028 23848 35080
rect 23900 35068 23906 35080
rect 24949 35071 25007 35077
rect 23900 35040 23945 35068
rect 23900 35028 23906 35040
rect 24949 35037 24961 35071
rect 24995 35064 25007 35071
rect 25038 35064 25044 35080
rect 24995 35037 25044 35064
rect 24949 35036 25044 35037
rect 24949 35031 25007 35036
rect 25038 35028 25044 35036
rect 25096 35028 25102 35080
rect 25682 35068 25688 35080
rect 25643 35040 25688 35068
rect 25682 35028 25688 35040
rect 25740 35028 25746 35080
rect 25869 35071 25927 35077
rect 25869 35037 25881 35071
rect 25915 35037 25927 35071
rect 25869 35031 25927 35037
rect 27065 35071 27123 35077
rect 27065 35037 27077 35071
rect 27111 35037 27123 35071
rect 27065 35031 27123 35037
rect 23106 35000 23112 35012
rect 22940 34972 23112 35000
rect 23106 34960 23112 34972
rect 23164 35000 23170 35012
rect 23474 35000 23480 35012
rect 23164 34972 23480 35000
rect 23164 34960 23170 34972
rect 23474 34960 23480 34972
rect 23532 35000 23538 35012
rect 25884 35000 25912 35031
rect 23532 34972 25912 35000
rect 27080 35000 27108 35031
rect 27522 35028 27528 35080
rect 27580 35068 27586 35080
rect 27985 35071 28043 35077
rect 27985 35068 27997 35071
rect 27580 35040 27997 35068
rect 27580 35028 27586 35040
rect 27985 35037 27997 35040
rect 28031 35037 28043 35071
rect 27985 35031 28043 35037
rect 28077 35071 28135 35077
rect 28077 35037 28089 35071
rect 28123 35037 28135 35071
rect 28077 35031 28135 35037
rect 27890 35000 27896 35012
rect 27080 34972 27896 35000
rect 23532 34960 23538 34972
rect 27890 34960 27896 34972
rect 27948 34960 27954 35012
rect 16945 34935 17003 34941
rect 16945 34901 16957 34935
rect 16991 34901 17003 34935
rect 16945 34895 17003 34901
rect 18601 34935 18659 34941
rect 18601 34901 18613 34935
rect 18647 34932 18659 34935
rect 19242 34932 19248 34944
rect 18647 34904 19248 34932
rect 18647 34901 18659 34904
rect 18601 34895 18659 34901
rect 19242 34892 19248 34904
rect 19300 34892 19306 34944
rect 22554 34892 22560 34944
rect 22612 34932 22618 34944
rect 23385 34935 23443 34941
rect 23385 34932 23397 34935
rect 22612 34904 23397 34932
rect 22612 34892 22618 34904
rect 23385 34901 23397 34904
rect 23431 34901 23443 34935
rect 23385 34895 23443 34901
rect 24854 34892 24860 34944
rect 24912 34932 24918 34944
rect 26050 34932 26056 34944
rect 24912 34904 26056 34932
rect 24912 34892 24918 34904
rect 26050 34892 26056 34904
rect 26108 34892 26114 34944
rect 26145 34935 26203 34941
rect 26145 34901 26157 34935
rect 26191 34932 26203 34935
rect 26326 34932 26332 34944
rect 26191 34904 26332 34932
rect 26191 34901 26203 34904
rect 26145 34895 26203 34901
rect 26326 34892 26332 34904
rect 26384 34932 26390 34944
rect 27430 34932 27436 34944
rect 26384 34904 27436 34932
rect 26384 34892 26390 34904
rect 27430 34892 27436 34904
rect 27488 34932 27494 34944
rect 28092 34932 28120 35031
rect 28166 35028 28172 35080
rect 28224 35068 28230 35080
rect 29914 35068 29920 35080
rect 28224 35040 28269 35068
rect 29875 35040 29920 35068
rect 28224 35028 28230 35040
rect 29914 35028 29920 35040
rect 29972 35028 29978 35080
rect 32030 35028 32036 35080
rect 32088 35068 32094 35080
rect 32769 35071 32827 35077
rect 32769 35068 32781 35071
rect 32088 35040 32781 35068
rect 32088 35028 32094 35040
rect 32769 35037 32781 35040
rect 32815 35068 32827 35071
rect 32858 35068 32864 35080
rect 32815 35040 32864 35068
rect 32815 35037 32827 35040
rect 32769 35031 32827 35037
rect 32858 35028 32864 35040
rect 32916 35068 32922 35080
rect 34701 35071 34759 35077
rect 34701 35068 34713 35071
rect 32916 35040 34713 35068
rect 32916 35028 32922 35040
rect 34701 35037 34713 35040
rect 34747 35068 34759 35071
rect 36170 35068 36176 35080
rect 34747 35040 36176 35068
rect 34747 35037 34759 35040
rect 34701 35031 34759 35037
rect 36170 35028 36176 35040
rect 36228 35028 36234 35080
rect 36725 35071 36783 35077
rect 36725 35037 36737 35071
rect 36771 35037 36783 35071
rect 37458 35068 37464 35080
rect 37419 35040 37464 35068
rect 36725 35031 36783 35037
rect 31846 35000 31852 35012
rect 31759 34972 31852 35000
rect 31846 34960 31852 34972
rect 31904 35000 31910 35012
rect 32122 35000 32128 35012
rect 31904 34972 32128 35000
rect 31904 34960 31910 34972
rect 32122 34960 32128 34972
rect 32180 34960 32186 35012
rect 33036 35003 33094 35009
rect 33036 34969 33048 35003
rect 33082 35000 33094 35003
rect 33226 35000 33232 35012
rect 33082 34972 33232 35000
rect 33082 34969 33094 34972
rect 33036 34963 33094 34969
rect 33226 34960 33232 34972
rect 33284 34960 33290 35012
rect 34790 34960 34796 35012
rect 34848 35000 34854 35012
rect 34946 35003 35004 35009
rect 34946 35000 34958 35003
rect 34848 34972 34958 35000
rect 34848 34960 34854 34972
rect 34946 34969 34958 34972
rect 34992 34969 35004 35003
rect 34946 34963 35004 34969
rect 35802 34960 35808 35012
rect 35860 35000 35866 35012
rect 36740 35000 36768 35031
rect 37458 35028 37464 35040
rect 37516 35028 37522 35080
rect 37553 35071 37611 35077
rect 37553 35037 37565 35071
rect 37599 35037 37611 35071
rect 37553 35031 37611 35037
rect 37568 35000 37596 35031
rect 35860 34972 37596 35000
rect 35860 34960 35866 34972
rect 27488 34904 28120 34932
rect 30193 34935 30251 34941
rect 27488 34892 27494 34904
rect 30193 34901 30205 34935
rect 30239 34932 30251 34935
rect 30466 34932 30472 34944
rect 30239 34904 30472 34932
rect 30239 34901 30251 34904
rect 30193 34895 30251 34901
rect 30466 34892 30472 34904
rect 30524 34892 30530 34944
rect 31938 34932 31944 34944
rect 31899 34904 31944 34932
rect 31938 34892 31944 34904
rect 31996 34892 32002 34944
rect 34149 34935 34207 34941
rect 34149 34901 34161 34935
rect 34195 34932 34207 34935
rect 34606 34932 34612 34944
rect 34195 34904 34612 34932
rect 34195 34901 34207 34904
rect 34149 34895 34207 34901
rect 34606 34892 34612 34904
rect 34664 34892 34670 34944
rect 37550 34892 37556 34944
rect 37608 34932 37614 34944
rect 37737 34935 37795 34941
rect 37737 34932 37749 34935
rect 37608 34904 37749 34932
rect 37608 34892 37614 34904
rect 37737 34901 37749 34904
rect 37783 34901 37795 34935
rect 37737 34895 37795 34901
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 15930 34728 15936 34740
rect 15891 34700 15936 34728
rect 15930 34688 15936 34700
rect 15988 34688 15994 34740
rect 18322 34728 18328 34740
rect 18283 34700 18328 34728
rect 18322 34688 18328 34700
rect 18380 34688 18386 34740
rect 20806 34728 20812 34740
rect 20767 34700 20812 34728
rect 20806 34688 20812 34700
rect 20864 34688 20870 34740
rect 22554 34688 22560 34740
rect 22612 34688 22618 34740
rect 23661 34731 23719 34737
rect 23661 34697 23673 34731
rect 23707 34728 23719 34731
rect 23842 34728 23848 34740
rect 23707 34700 23848 34728
rect 23707 34697 23719 34700
rect 23661 34691 23719 34697
rect 23842 34688 23848 34700
rect 23900 34688 23906 34740
rect 26970 34728 26976 34740
rect 23952 34700 26976 34728
rect 17218 34669 17224 34672
rect 17212 34660 17224 34669
rect 17179 34632 17224 34660
rect 17212 34623 17224 34632
rect 17218 34620 17224 34623
rect 17276 34620 17282 34672
rect 22563 34607 22591 34688
rect 22830 34660 22836 34672
rect 22667 34632 22836 34660
rect 16117 34595 16175 34601
rect 16117 34561 16129 34595
rect 16163 34592 16175 34595
rect 16666 34592 16672 34604
rect 16163 34564 16672 34592
rect 16163 34561 16175 34564
rect 16117 34555 16175 34561
rect 16666 34552 16672 34564
rect 16724 34552 16730 34604
rect 19426 34552 19432 34604
rect 19484 34592 19490 34604
rect 19898 34595 19956 34601
rect 19898 34592 19910 34595
rect 19484 34564 19910 34592
rect 19484 34552 19490 34564
rect 19898 34561 19910 34564
rect 19944 34561 19956 34595
rect 19898 34555 19956 34561
rect 20993 34595 21051 34601
rect 20993 34561 21005 34595
rect 21039 34592 21051 34595
rect 21082 34592 21088 34604
rect 21039 34564 21088 34592
rect 21039 34561 21051 34564
rect 20993 34555 21051 34561
rect 21082 34552 21088 34564
rect 21140 34552 21146 34604
rect 21177 34595 21235 34601
rect 21177 34561 21189 34595
rect 21223 34592 21235 34595
rect 21266 34592 21272 34604
rect 21223 34564 21272 34592
rect 21223 34561 21235 34564
rect 21177 34555 21235 34561
rect 21266 34552 21272 34564
rect 21324 34552 21330 34604
rect 21634 34552 21640 34604
rect 21692 34592 21698 34604
rect 22552 34601 22610 34607
rect 22667 34604 22695 34632
rect 22830 34620 22836 34632
rect 22888 34660 22894 34672
rect 23952 34660 23980 34700
rect 26970 34688 26976 34700
rect 27028 34688 27034 34740
rect 29914 34728 29920 34740
rect 29196 34700 29920 34728
rect 26326 34660 26332 34672
rect 22888 34632 23980 34660
rect 26252 34632 26332 34660
rect 22888 34620 22894 34632
rect 22373 34595 22431 34601
rect 22373 34592 22385 34595
rect 21692 34564 22385 34592
rect 21692 34552 21698 34564
rect 22373 34561 22385 34564
rect 22419 34561 22431 34595
rect 22552 34567 22564 34601
rect 22598 34567 22610 34601
rect 22552 34561 22610 34567
rect 22652 34598 22710 34604
rect 22652 34564 22664 34598
rect 22698 34564 22710 34598
rect 22373 34555 22431 34561
rect 22652 34558 22710 34564
rect 22738 34552 22744 34604
rect 22796 34592 22802 34604
rect 23474 34592 23480 34604
rect 22796 34564 23336 34592
rect 23435 34564 23480 34592
rect 22796 34552 22802 34564
rect 15194 34484 15200 34536
rect 15252 34524 15258 34536
rect 15562 34524 15568 34536
rect 15252 34496 15568 34524
rect 15252 34484 15258 34496
rect 15562 34484 15568 34496
rect 15620 34524 15626 34536
rect 16482 34524 16488 34536
rect 15620 34496 16488 34524
rect 15620 34484 15626 34496
rect 16482 34484 16488 34496
rect 16540 34524 16546 34536
rect 16945 34527 17003 34533
rect 16945 34524 16957 34527
rect 16540 34496 16957 34524
rect 16540 34484 16546 34496
rect 16945 34493 16957 34496
rect 16991 34493 17003 34527
rect 20162 34524 20168 34536
rect 20123 34496 20168 34524
rect 16945 34487 17003 34493
rect 20162 34484 20168 34496
rect 20220 34484 20226 34536
rect 22830 34484 22836 34536
rect 22888 34524 22894 34536
rect 23017 34527 23075 34533
rect 23017 34524 23029 34527
rect 22888 34496 23029 34524
rect 22888 34484 22894 34496
rect 23017 34493 23029 34496
rect 23063 34493 23075 34527
rect 23308 34524 23336 34564
rect 23474 34552 23480 34564
rect 23532 34552 23538 34604
rect 23566 34552 23572 34604
rect 23624 34592 23630 34604
rect 23661 34595 23719 34601
rect 23661 34592 23673 34595
rect 23624 34564 23673 34592
rect 23624 34552 23630 34564
rect 23661 34561 23673 34564
rect 23707 34561 23719 34595
rect 23661 34555 23719 34561
rect 24302 34552 24308 34604
rect 24360 34592 24366 34604
rect 24489 34595 24547 34601
rect 24489 34592 24501 34595
rect 24360 34564 24501 34592
rect 24360 34552 24366 34564
rect 24489 34561 24501 34564
rect 24535 34561 24547 34595
rect 24670 34592 24676 34604
rect 24631 34564 24676 34592
rect 24489 34555 24547 34561
rect 24670 34552 24676 34564
rect 24728 34552 24734 34604
rect 24762 34552 24768 34604
rect 24820 34592 24826 34604
rect 25038 34592 25044 34604
rect 24820 34564 24865 34592
rect 24951 34564 25044 34592
rect 24820 34552 24826 34564
rect 25038 34552 25044 34564
rect 25096 34592 25102 34604
rect 26252 34601 26280 34632
rect 26326 34620 26332 34632
rect 26384 34620 26390 34672
rect 26237 34595 26295 34601
rect 25096 34564 25636 34592
rect 25096 34552 25102 34564
rect 24854 34524 24860 34536
rect 23308 34496 24532 34524
rect 24815 34496 24860 34524
rect 23017 34487 23075 34493
rect 24504 34468 24532 34496
rect 24854 34484 24860 34496
rect 24912 34484 24918 34536
rect 24486 34416 24492 34468
rect 24544 34416 24550 34468
rect 25608 34456 25636 34564
rect 26237 34561 26249 34595
rect 26283 34561 26295 34595
rect 26418 34592 26424 34604
rect 26379 34564 26424 34592
rect 26237 34555 26295 34561
rect 26418 34552 26424 34564
rect 26476 34552 26482 34604
rect 26602 34552 26608 34604
rect 26660 34592 26666 34604
rect 27157 34595 27215 34601
rect 27157 34592 27169 34595
rect 26660 34564 27169 34592
rect 26660 34552 26666 34564
rect 27157 34561 27169 34564
rect 27203 34561 27215 34595
rect 27338 34592 27344 34604
rect 27299 34564 27344 34592
rect 27157 34555 27215 34561
rect 27338 34552 27344 34564
rect 27396 34552 27402 34604
rect 27433 34595 27491 34601
rect 27433 34561 27445 34595
rect 27479 34561 27491 34595
rect 27433 34555 27491 34561
rect 26329 34527 26387 34533
rect 26329 34493 26341 34527
rect 26375 34524 26387 34527
rect 27448 34524 27476 34555
rect 27706 34552 27712 34604
rect 27764 34592 27770 34604
rect 28353 34595 28411 34601
rect 28353 34592 28365 34595
rect 27764 34564 28365 34592
rect 27764 34552 27770 34564
rect 28353 34561 28365 34564
rect 28399 34561 28411 34595
rect 28353 34555 28411 34561
rect 28442 34552 28448 34604
rect 28500 34592 28506 34604
rect 29196 34601 29224 34700
rect 29914 34688 29920 34700
rect 29972 34728 29978 34740
rect 30009 34731 30067 34737
rect 30009 34728 30021 34731
rect 29972 34700 30021 34728
rect 29972 34688 29978 34700
rect 30009 34697 30021 34700
rect 30055 34697 30067 34731
rect 30009 34691 30067 34697
rect 33226 34688 33232 34740
rect 33284 34728 33290 34740
rect 33505 34731 33563 34737
rect 33505 34728 33517 34731
rect 33284 34700 33517 34728
rect 33284 34688 33290 34700
rect 33505 34697 33517 34700
rect 33551 34697 33563 34731
rect 33505 34691 33563 34697
rect 34514 34688 34520 34740
rect 34572 34728 34578 34740
rect 36173 34731 36231 34737
rect 36173 34728 36185 34731
rect 34572 34700 36185 34728
rect 34572 34688 34578 34700
rect 36173 34697 36185 34700
rect 36219 34697 36231 34731
rect 36173 34691 36231 34697
rect 36998 34688 37004 34740
rect 37056 34728 37062 34740
rect 37369 34731 37427 34737
rect 37369 34728 37381 34731
rect 37056 34700 37381 34728
rect 37056 34688 37062 34700
rect 37369 34697 37381 34700
rect 37415 34697 37427 34731
rect 37369 34691 37427 34697
rect 32392 34663 32450 34669
rect 32392 34629 32404 34663
rect 32438 34660 32450 34663
rect 32582 34660 32588 34672
rect 32438 34632 32588 34660
rect 32438 34629 32450 34632
rect 32392 34623 32450 34629
rect 32582 34620 32588 34632
rect 32640 34620 32646 34672
rect 34606 34620 34612 34672
rect 34664 34660 34670 34672
rect 35713 34663 35771 34669
rect 35713 34660 35725 34663
rect 34664 34632 35725 34660
rect 34664 34620 34670 34632
rect 35713 34629 35725 34632
rect 35759 34629 35771 34663
rect 35713 34623 35771 34629
rect 35894 34620 35900 34672
rect 35952 34660 35958 34672
rect 36325 34663 36383 34669
rect 36325 34660 36337 34663
rect 35952 34632 36337 34660
rect 35952 34620 35958 34632
rect 36325 34629 36337 34632
rect 36371 34629 36383 34663
rect 36325 34623 36383 34629
rect 36541 34663 36599 34669
rect 36541 34629 36553 34663
rect 36587 34660 36599 34663
rect 36722 34660 36728 34672
rect 36587 34632 36728 34660
rect 36587 34629 36599 34632
rect 36541 34623 36599 34629
rect 29181 34595 29239 34601
rect 29181 34592 29193 34595
rect 28500 34564 29193 34592
rect 28500 34552 28506 34564
rect 29181 34561 29193 34564
rect 29227 34561 29239 34595
rect 29181 34555 29239 34561
rect 30558 34552 30564 34604
rect 30616 34592 30622 34604
rect 31122 34595 31180 34601
rect 31122 34592 31134 34595
rect 30616 34564 31134 34592
rect 30616 34552 30622 34564
rect 31122 34561 31134 34564
rect 31168 34561 31180 34595
rect 31122 34555 31180 34561
rect 34241 34595 34299 34601
rect 34241 34561 34253 34595
rect 34287 34592 34299 34595
rect 34422 34592 34428 34604
rect 34287 34564 34428 34592
rect 34287 34561 34299 34564
rect 34241 34555 34299 34561
rect 34422 34552 34428 34564
rect 34480 34552 34486 34604
rect 35434 34592 35440 34604
rect 35395 34564 35440 34592
rect 35434 34552 35440 34564
rect 35492 34552 35498 34604
rect 27893 34527 27951 34533
rect 27893 34524 27905 34527
rect 26375 34496 27905 34524
rect 26375 34493 26387 34496
rect 26329 34487 26387 34493
rect 27893 34493 27905 34496
rect 27939 34493 27951 34527
rect 27893 34487 27951 34493
rect 27982 34484 27988 34536
rect 28040 34524 28046 34536
rect 28258 34524 28264 34536
rect 28040 34496 28264 34524
rect 28040 34484 28046 34496
rect 28258 34484 28264 34496
rect 28316 34484 28322 34536
rect 28537 34527 28595 34533
rect 28537 34493 28549 34527
rect 28583 34524 28595 34527
rect 29086 34524 29092 34536
rect 28583 34496 29092 34524
rect 28583 34493 28595 34496
rect 28537 34487 28595 34493
rect 29086 34484 29092 34496
rect 29144 34484 29150 34536
rect 29273 34527 29331 34533
rect 29273 34524 29285 34527
rect 29196 34496 29285 34524
rect 26418 34456 26424 34468
rect 25608 34428 26424 34456
rect 26418 34416 26424 34428
rect 26476 34416 26482 34468
rect 28074 34416 28080 34468
rect 28132 34456 28138 34468
rect 29196 34456 29224 34496
rect 29273 34493 29285 34496
rect 29319 34493 29331 34527
rect 29546 34524 29552 34536
rect 29507 34496 29552 34524
rect 29273 34487 29331 34493
rect 29546 34484 29552 34496
rect 29604 34484 29610 34536
rect 31389 34527 31447 34533
rect 31389 34493 31401 34527
rect 31435 34524 31447 34527
rect 32030 34524 32036 34536
rect 31435 34496 32036 34524
rect 31435 34493 31447 34496
rect 31389 34487 31447 34493
rect 32030 34484 32036 34496
rect 32088 34524 32094 34536
rect 32125 34527 32183 34533
rect 32125 34524 32137 34527
rect 32088 34496 32137 34524
rect 32088 34484 32094 34496
rect 32125 34493 32137 34496
rect 32171 34493 32183 34527
rect 33962 34524 33968 34536
rect 33923 34496 33968 34524
rect 32125 34487 32183 34493
rect 33962 34484 33968 34496
rect 34020 34484 34026 34536
rect 35621 34527 35679 34533
rect 35621 34493 35633 34527
rect 35667 34524 35679 34527
rect 36354 34524 36360 34536
rect 35667 34496 36360 34524
rect 35667 34493 35679 34496
rect 35621 34487 35679 34493
rect 36354 34484 36360 34496
rect 36412 34484 36418 34536
rect 36556 34456 36584 34623
rect 36722 34620 36728 34632
rect 36780 34620 36786 34672
rect 37550 34592 37556 34604
rect 37511 34564 37556 34592
rect 37550 34552 37556 34564
rect 37608 34552 37614 34604
rect 28132 34428 29224 34456
rect 35728 34428 36584 34456
rect 28132 34416 28138 34428
rect 18138 34348 18144 34400
rect 18196 34388 18202 34400
rect 18785 34391 18843 34397
rect 18785 34388 18797 34391
rect 18196 34360 18797 34388
rect 18196 34348 18202 34360
rect 18785 34357 18797 34360
rect 18831 34357 18843 34391
rect 18785 34351 18843 34357
rect 25225 34391 25283 34397
rect 25225 34357 25237 34391
rect 25271 34388 25283 34391
rect 25314 34388 25320 34400
rect 25271 34360 25320 34388
rect 25271 34357 25283 34360
rect 25225 34351 25283 34357
rect 25314 34348 25320 34360
rect 25372 34348 25378 34400
rect 26878 34348 26884 34400
rect 26936 34388 26942 34400
rect 26973 34391 27031 34397
rect 26973 34388 26985 34391
rect 26936 34360 26985 34388
rect 26936 34348 26942 34360
rect 26973 34357 26985 34360
rect 27019 34357 27031 34391
rect 26973 34351 27031 34357
rect 34790 34348 34796 34400
rect 34848 34388 34854 34400
rect 35728 34397 35756 34428
rect 35253 34391 35311 34397
rect 35253 34388 35265 34391
rect 34848 34360 35265 34388
rect 34848 34348 34854 34360
rect 35253 34357 35265 34360
rect 35299 34357 35311 34391
rect 35253 34351 35311 34357
rect 35713 34391 35771 34397
rect 35713 34357 35725 34391
rect 35759 34357 35771 34391
rect 36354 34388 36360 34400
rect 36315 34360 36360 34388
rect 35713 34351 35771 34357
rect 36354 34348 36360 34360
rect 36412 34348 36418 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 16666 34184 16672 34196
rect 16627 34156 16672 34184
rect 16666 34144 16672 34156
rect 16724 34144 16730 34196
rect 19426 34184 19432 34196
rect 19387 34156 19432 34184
rect 19426 34144 19432 34156
rect 19484 34144 19490 34196
rect 24857 34187 24915 34193
rect 24857 34153 24869 34187
rect 24903 34184 24915 34187
rect 25682 34184 25688 34196
rect 24903 34156 25688 34184
rect 24903 34153 24915 34156
rect 24857 34147 24915 34153
rect 25682 34144 25688 34156
rect 25740 34144 25746 34196
rect 27893 34187 27951 34193
rect 27893 34153 27905 34187
rect 27939 34184 27951 34187
rect 28166 34184 28172 34196
rect 27939 34156 28172 34184
rect 27939 34153 27951 34156
rect 27893 34147 27951 34153
rect 28166 34144 28172 34156
rect 28224 34144 28230 34196
rect 30558 34184 30564 34196
rect 30519 34156 30564 34184
rect 30558 34144 30564 34156
rect 30616 34144 30622 34196
rect 34698 34184 34704 34196
rect 34659 34156 34704 34184
rect 34698 34144 34704 34156
rect 34756 34144 34762 34196
rect 35713 34187 35771 34193
rect 35713 34153 35725 34187
rect 35759 34184 35771 34187
rect 35894 34184 35900 34196
rect 35759 34156 35900 34184
rect 35759 34153 35771 34156
rect 35713 34147 35771 34153
rect 35894 34144 35900 34156
rect 35952 34144 35958 34196
rect 37734 34184 37740 34196
rect 36740 34156 37740 34184
rect 16209 34119 16267 34125
rect 16209 34085 16221 34119
rect 16255 34116 16267 34119
rect 17862 34116 17868 34128
rect 16255 34088 16574 34116
rect 17823 34088 17868 34116
rect 16255 34085 16267 34088
rect 16209 34079 16267 34085
rect 16546 34048 16574 34088
rect 17862 34076 17868 34088
rect 17920 34076 17926 34128
rect 30101 34119 30159 34125
rect 30101 34085 30113 34119
rect 30147 34085 30159 34119
rect 30101 34079 30159 34085
rect 24397 34051 24455 34057
rect 16546 34020 17080 34048
rect 14829 33983 14887 33989
rect 14829 33949 14841 33983
rect 14875 33980 14887 33983
rect 16850 33980 16856 33992
rect 14875 33952 15240 33980
rect 16811 33952 16856 33980
rect 14875 33949 14887 33952
rect 14829 33943 14887 33949
rect 15212 33924 15240 33952
rect 16850 33940 16856 33952
rect 16908 33940 16914 33992
rect 17052 33989 17080 34020
rect 24397 34017 24409 34051
rect 24443 34048 24455 34051
rect 25038 34048 25044 34060
rect 24443 34020 25044 34048
rect 24443 34017 24455 34020
rect 24397 34011 24455 34017
rect 25038 34008 25044 34020
rect 25096 34008 25102 34060
rect 26786 34048 26792 34060
rect 26699 34020 26792 34048
rect 17037 33983 17095 33989
rect 17037 33949 17049 33983
rect 17083 33949 17095 33983
rect 18138 33980 18144 33992
rect 18099 33952 18144 33980
rect 17037 33943 17095 33949
rect 15102 33921 15108 33924
rect 15096 33912 15108 33921
rect 15063 33884 15108 33912
rect 15096 33875 15108 33884
rect 15102 33872 15108 33875
rect 15160 33872 15166 33924
rect 15194 33872 15200 33924
rect 15252 33872 15258 33924
rect 17052 33912 17080 33943
rect 18138 33940 18144 33952
rect 18196 33940 18202 33992
rect 18233 33983 18291 33989
rect 18233 33949 18245 33983
rect 18279 33980 18291 33983
rect 18322 33980 18328 33992
rect 18279 33952 18328 33980
rect 18279 33949 18291 33952
rect 18233 33943 18291 33949
rect 18322 33940 18328 33952
rect 18380 33940 18386 33992
rect 19242 33980 19248 33992
rect 19203 33952 19248 33980
rect 19242 33940 19248 33952
rect 19300 33940 19306 33992
rect 20162 33940 20168 33992
rect 20220 33980 20226 33992
rect 21361 33983 21419 33989
rect 21361 33980 21373 33983
rect 20220 33952 21373 33980
rect 20220 33940 20226 33952
rect 21361 33949 21373 33952
rect 21407 33980 21419 33983
rect 23014 33980 23020 33992
rect 21407 33952 23020 33980
rect 21407 33949 21419 33952
rect 21361 33943 21419 33949
rect 23014 33940 23020 33952
rect 23072 33940 23078 33992
rect 24486 33980 24492 33992
rect 24447 33952 24492 33980
rect 24486 33940 24492 33952
rect 24544 33940 24550 33992
rect 24673 33983 24731 33989
rect 24673 33949 24685 33983
rect 24719 33980 24731 33983
rect 24946 33980 24952 33992
rect 24719 33952 24952 33980
rect 24719 33949 24731 33952
rect 24673 33943 24731 33949
rect 24946 33940 24952 33952
rect 25004 33940 25010 33992
rect 26712 33989 26740 34020
rect 26786 34008 26792 34020
rect 26844 34048 26850 34060
rect 26844 34020 28580 34048
rect 26844 34008 26850 34020
rect 26697 33983 26755 33989
rect 26697 33949 26709 33983
rect 26743 33949 26755 33983
rect 26878 33980 26884 33992
rect 26839 33952 26884 33980
rect 26697 33943 26755 33949
rect 26878 33940 26884 33952
rect 26936 33940 26942 33992
rect 26970 33940 26976 33992
rect 27028 33980 27034 33992
rect 27111 33983 27169 33989
rect 27028 33952 27073 33980
rect 27028 33940 27034 33952
rect 27111 33949 27123 33983
rect 27157 33980 27169 33983
rect 28074 33980 28080 33992
rect 27157 33952 27936 33980
rect 28035 33952 28080 33980
rect 27157 33949 27169 33952
rect 27111 33943 27169 33949
rect 17052 33884 18092 33912
rect 18064 33856 18092 33884
rect 20898 33872 20904 33924
rect 20956 33912 20962 33924
rect 21094 33915 21152 33921
rect 21094 33912 21106 33915
rect 20956 33884 21106 33912
rect 20956 33872 20962 33884
rect 21094 33881 21106 33884
rect 21140 33881 21152 33915
rect 27908 33912 27936 33952
rect 28074 33940 28080 33952
rect 28132 33940 28138 33992
rect 28258 33980 28264 33992
rect 28219 33952 28264 33980
rect 28258 33940 28264 33952
rect 28316 33940 28322 33992
rect 28353 33983 28411 33989
rect 28353 33949 28365 33983
rect 28399 33980 28411 33983
rect 28442 33980 28448 33992
rect 28399 33952 28448 33980
rect 28399 33949 28411 33952
rect 28353 33943 28411 33949
rect 28442 33940 28448 33952
rect 28500 33940 28506 33992
rect 28276 33912 28304 33940
rect 27908 33884 28304 33912
rect 28552 33912 28580 34020
rect 29086 34008 29092 34060
rect 29144 34048 29150 34060
rect 29641 34051 29699 34057
rect 29641 34048 29653 34051
rect 29144 34020 29653 34048
rect 29144 34008 29150 34020
rect 29641 34017 29653 34020
rect 29687 34017 29699 34051
rect 30116 34048 30144 34079
rect 30650 34076 30656 34128
rect 30708 34116 30714 34128
rect 32950 34116 32956 34128
rect 30708 34088 32956 34116
rect 30708 34076 30714 34088
rect 32950 34076 32956 34088
rect 33008 34116 33014 34128
rect 36740 34116 36768 34156
rect 37734 34144 37740 34156
rect 37792 34144 37798 34196
rect 33008 34088 34100 34116
rect 33008 34076 33014 34088
rect 32122 34048 32128 34060
rect 30116 34020 30880 34048
rect 32083 34020 32128 34048
rect 29641 34011 29699 34017
rect 29546 33940 29552 33992
rect 29604 33980 29610 33992
rect 29733 33983 29791 33989
rect 29733 33980 29745 33983
rect 29604 33952 29745 33980
rect 29604 33940 29610 33952
rect 29733 33949 29745 33952
rect 29779 33949 29791 33983
rect 29733 33943 29791 33949
rect 30466 33940 30472 33992
rect 30524 33980 30530 33992
rect 30852 33989 30880 34020
rect 32122 34008 32128 34020
rect 32180 34008 32186 34060
rect 33778 34048 33784 34060
rect 33739 34020 33784 34048
rect 33778 34008 33784 34020
rect 33836 34008 33842 34060
rect 34072 34057 34100 34088
rect 35912 34088 36768 34116
rect 34057 34051 34115 34057
rect 34057 34017 34069 34051
rect 34103 34017 34115 34051
rect 34057 34011 34115 34017
rect 34149 34051 34207 34057
rect 34149 34017 34161 34051
rect 34195 34048 34207 34051
rect 34514 34048 34520 34060
rect 34195 34020 34520 34048
rect 34195 34017 34207 34020
rect 34149 34011 34207 34017
rect 34514 34008 34520 34020
rect 34572 34008 34578 34060
rect 35802 34048 35808 34060
rect 34900 34020 35808 34048
rect 30561 33983 30619 33989
rect 30561 33980 30573 33983
rect 30524 33952 30573 33980
rect 30524 33940 30530 33952
rect 30561 33949 30573 33952
rect 30607 33949 30619 33983
rect 30561 33943 30619 33949
rect 30837 33983 30895 33989
rect 30837 33949 30849 33983
rect 30883 33949 30895 33983
rect 30837 33943 30895 33949
rect 32214 33940 32220 33992
rect 32272 33980 32278 33992
rect 32401 33983 32459 33989
rect 32401 33980 32413 33983
rect 32272 33952 32413 33980
rect 32272 33940 32278 33952
rect 32401 33949 32413 33952
rect 32447 33949 32459 33983
rect 33686 33980 33692 33992
rect 33647 33952 33692 33980
rect 32401 33943 32459 33949
rect 33686 33940 33692 33952
rect 33744 33940 33750 33992
rect 34900 33989 34928 34020
rect 35802 34008 35808 34020
rect 35860 34008 35866 34060
rect 35912 33989 35940 34088
rect 36170 34008 36176 34060
rect 36228 34048 36234 34060
rect 36725 34051 36783 34057
rect 36725 34048 36737 34051
rect 36228 34020 36737 34048
rect 36228 34008 36234 34020
rect 36725 34017 36737 34020
rect 36771 34017 36783 34051
rect 36725 34011 36783 34017
rect 34885 33983 34943 33989
rect 34885 33949 34897 33983
rect 34931 33949 34943 33983
rect 34885 33943 34943 33949
rect 34977 33983 35035 33989
rect 34977 33949 34989 33983
rect 35023 33949 35035 33983
rect 34977 33943 35035 33949
rect 35897 33983 35955 33989
rect 35897 33949 35909 33983
rect 35943 33949 35955 33983
rect 35897 33943 35955 33949
rect 36081 33983 36139 33989
rect 36081 33949 36093 33983
rect 36127 33980 36139 33983
rect 37458 33980 37464 33992
rect 36127 33952 37464 33980
rect 36127 33949 36139 33952
rect 36081 33943 36139 33949
rect 34606 33912 34612 33924
rect 28552 33884 31754 33912
rect 21094 33875 21152 33881
rect 18046 33844 18052 33856
rect 18007 33816 18052 33844
rect 18046 33804 18052 33816
rect 18104 33804 18110 33856
rect 18414 33844 18420 33856
rect 18375 33816 18420 33844
rect 18414 33804 18420 33816
rect 18472 33804 18478 33856
rect 19981 33847 20039 33853
rect 19981 33813 19993 33847
rect 20027 33844 20039 33847
rect 20070 33844 20076 33856
rect 20027 33816 20076 33844
rect 20027 33813 20039 33816
rect 19981 33807 20039 33813
rect 20070 33804 20076 33816
rect 20128 33804 20134 33856
rect 27341 33847 27399 33853
rect 27341 33813 27353 33847
rect 27387 33844 27399 33847
rect 28534 33844 28540 33856
rect 27387 33816 28540 33844
rect 27387 33813 27399 33816
rect 27341 33807 27399 33813
rect 28534 33804 28540 33816
rect 28592 33804 28598 33856
rect 29822 33804 29828 33856
rect 29880 33844 29886 33856
rect 30745 33847 30803 33853
rect 30745 33844 30757 33847
rect 29880 33816 30757 33844
rect 29880 33804 29886 33816
rect 30745 33813 30757 33816
rect 30791 33813 30803 33847
rect 31726 33844 31754 33884
rect 33980 33884 34612 33912
rect 31938 33844 31944 33856
rect 31726 33816 31944 33844
rect 30745 33807 30803 33813
rect 31938 33804 31944 33816
rect 31996 33844 32002 33856
rect 33318 33844 33324 33856
rect 31996 33816 33324 33844
rect 31996 33804 32002 33816
rect 33318 33804 33324 33816
rect 33376 33804 33382 33856
rect 33502 33844 33508 33856
rect 33463 33816 33508 33844
rect 33502 33804 33508 33816
rect 33560 33804 33566 33856
rect 33980 33853 34008 33884
rect 34606 33872 34612 33884
rect 34664 33912 34670 33924
rect 34992 33912 35020 33943
rect 37458 33940 37464 33952
rect 37516 33940 37522 33992
rect 34664 33884 35020 33912
rect 35989 33915 36047 33921
rect 34664 33872 34670 33884
rect 35989 33881 36001 33915
rect 36035 33912 36047 33915
rect 36035 33884 36216 33912
rect 36035 33881 36047 33884
rect 35989 33875 36047 33881
rect 33965 33847 34023 33853
rect 33965 33813 33977 33847
rect 34011 33813 34023 33847
rect 36188 33844 36216 33884
rect 36262 33872 36268 33924
rect 36320 33912 36326 33924
rect 36998 33921 37004 33924
rect 36320 33884 36365 33912
rect 36320 33872 36326 33884
rect 36992 33875 37004 33921
rect 37056 33912 37062 33924
rect 37056 33884 37092 33912
rect 36998 33872 37004 33875
rect 37056 33872 37062 33884
rect 37550 33844 37556 33856
rect 36188 33816 37556 33844
rect 33965 33807 34023 33813
rect 37550 33804 37556 33816
rect 37608 33804 37614 33856
rect 38102 33844 38108 33856
rect 38063 33816 38108 33844
rect 38102 33804 38108 33816
rect 38160 33804 38166 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 15102 33600 15108 33652
rect 15160 33640 15166 33652
rect 15197 33643 15255 33649
rect 15197 33640 15209 33643
rect 15160 33612 15209 33640
rect 15160 33600 15166 33612
rect 15197 33609 15209 33612
rect 15243 33609 15255 33643
rect 15197 33603 15255 33609
rect 17773 33643 17831 33649
rect 17773 33609 17785 33643
rect 17819 33640 17831 33643
rect 17954 33640 17960 33652
rect 17819 33612 17960 33640
rect 17819 33609 17831 33612
rect 17773 33603 17831 33609
rect 17954 33600 17960 33612
rect 18012 33600 18018 33652
rect 27157 33643 27215 33649
rect 27157 33609 27169 33643
rect 27203 33640 27215 33643
rect 27338 33640 27344 33652
rect 27203 33612 27344 33640
rect 27203 33609 27215 33612
rect 27157 33603 27215 33609
rect 27338 33600 27344 33612
rect 27396 33600 27402 33652
rect 30561 33643 30619 33649
rect 30561 33609 30573 33643
rect 30607 33640 30619 33643
rect 30650 33640 30656 33652
rect 30607 33612 30656 33640
rect 30607 33609 30619 33612
rect 30561 33603 30619 33609
rect 30650 33600 30656 33612
rect 30708 33600 30714 33652
rect 33686 33600 33692 33652
rect 33744 33640 33750 33652
rect 34241 33643 34299 33649
rect 34241 33640 34253 33643
rect 33744 33612 34253 33640
rect 33744 33600 33750 33612
rect 34241 33609 34253 33612
rect 34287 33609 34299 33643
rect 34241 33603 34299 33609
rect 18233 33575 18291 33581
rect 18233 33541 18245 33575
rect 18279 33572 18291 33575
rect 18322 33572 18328 33584
rect 18279 33544 18328 33572
rect 18279 33541 18291 33544
rect 18233 33535 18291 33541
rect 18322 33532 18328 33544
rect 18380 33532 18386 33584
rect 21082 33532 21088 33584
rect 21140 33572 21146 33584
rect 27522 33572 27528 33584
rect 21140 33544 27200 33572
rect 27483 33544 27528 33572
rect 21140 33532 21146 33544
rect 15378 33504 15384 33516
rect 15339 33476 15384 33504
rect 15378 33464 15384 33476
rect 15436 33464 15442 33516
rect 17862 33464 17868 33516
rect 17920 33504 17926 33516
rect 17957 33507 18015 33513
rect 17957 33504 17969 33507
rect 17920 33476 17969 33504
rect 17920 33464 17926 33476
rect 17957 33473 17969 33476
rect 18003 33473 18015 33507
rect 20990 33504 20996 33516
rect 20951 33476 20996 33504
rect 17957 33467 18015 33473
rect 20990 33464 20996 33476
rect 21048 33464 21054 33516
rect 21836 33513 21864 33544
rect 21821 33507 21879 33513
rect 21821 33473 21833 33507
rect 21867 33473 21879 33507
rect 21821 33467 21879 33473
rect 23014 33464 23020 33516
rect 23072 33504 23078 33516
rect 25314 33513 25320 33516
rect 25041 33507 25099 33513
rect 25041 33504 25053 33507
rect 23072 33476 25053 33504
rect 23072 33464 23078 33476
rect 25041 33473 25053 33476
rect 25087 33473 25099 33507
rect 25308 33504 25320 33513
rect 25275 33476 25320 33504
rect 25041 33467 25099 33473
rect 25308 33467 25320 33476
rect 25314 33464 25320 33467
rect 25372 33464 25378 33516
rect 18138 33436 18144 33448
rect 18099 33408 18144 33436
rect 18138 33396 18144 33408
rect 18196 33396 18202 33448
rect 27172 33436 27200 33544
rect 27522 33532 27528 33544
rect 27580 33532 27586 33584
rect 29638 33572 29644 33584
rect 29599 33544 29644 33572
rect 29638 33532 29644 33544
rect 29696 33532 29702 33584
rect 36262 33532 36268 33584
rect 36320 33572 36326 33584
rect 38102 33572 38108 33584
rect 36320 33544 38108 33572
rect 36320 33532 36326 33544
rect 27341 33507 27399 33513
rect 27341 33473 27353 33507
rect 27387 33504 27399 33507
rect 27430 33504 27436 33516
rect 27387 33476 27436 33504
rect 27387 33473 27399 33476
rect 27341 33467 27399 33473
rect 27430 33464 27436 33476
rect 27488 33464 27494 33516
rect 30374 33504 30380 33516
rect 30335 33476 30380 33504
rect 30374 33464 30380 33476
rect 30432 33464 30438 33516
rect 34422 33504 34428 33516
rect 34383 33476 34428 33504
rect 34422 33464 34428 33476
rect 34480 33464 34486 33516
rect 34701 33507 34759 33513
rect 34701 33473 34713 33507
rect 34747 33504 34759 33507
rect 34790 33504 34796 33516
rect 34747 33476 34796 33504
rect 34747 33473 34759 33476
rect 34701 33467 34759 33473
rect 34790 33464 34796 33476
rect 34848 33464 34854 33516
rect 36633 33507 36691 33513
rect 36633 33473 36645 33507
rect 36679 33504 36691 33507
rect 37274 33504 37280 33516
rect 36679 33476 37280 33504
rect 36679 33473 36691 33476
rect 36633 33467 36691 33473
rect 37274 33464 37280 33476
rect 37332 33464 37338 33516
rect 37476 33513 37504 33544
rect 38102 33532 38108 33544
rect 38160 33532 38166 33584
rect 37461 33507 37519 33513
rect 37461 33473 37473 33507
rect 37507 33473 37519 33507
rect 37461 33467 37519 33473
rect 37550 33464 37556 33516
rect 37608 33504 37614 33516
rect 37608 33476 37653 33504
rect 37608 33464 37614 33476
rect 37734 33464 37740 33516
rect 37792 33504 37798 33516
rect 37792 33476 37837 33504
rect 37792 33464 37798 33476
rect 31294 33436 31300 33448
rect 27172 33408 31300 33436
rect 31294 33396 31300 33408
rect 31352 33396 31358 33448
rect 21177 33371 21235 33377
rect 21177 33337 21189 33371
rect 21223 33368 21235 33371
rect 21818 33368 21824 33380
rect 21223 33340 21824 33368
rect 21223 33337 21235 33340
rect 21177 33331 21235 33337
rect 21818 33328 21824 33340
rect 21876 33368 21882 33380
rect 23106 33368 23112 33380
rect 21876 33340 23112 33368
rect 21876 33328 21882 33340
rect 23106 33328 23112 33340
rect 23164 33328 23170 33380
rect 33962 33368 33968 33380
rect 25976 33340 33968 33368
rect 18046 33300 18052 33312
rect 18007 33272 18052 33300
rect 18046 33260 18052 33272
rect 18104 33260 18110 33312
rect 22002 33300 22008 33312
rect 21915 33272 22008 33300
rect 22002 33260 22008 33272
rect 22060 33300 22066 33312
rect 22830 33300 22836 33312
rect 22060 33272 22836 33300
rect 22060 33260 22066 33272
rect 22830 33260 22836 33272
rect 22888 33300 22894 33312
rect 25976 33300 26004 33340
rect 33962 33328 33968 33340
rect 34020 33368 34026 33380
rect 34514 33368 34520 33380
rect 34020 33340 34520 33368
rect 34020 33328 34026 33340
rect 34514 33328 34520 33340
rect 34572 33328 34578 33380
rect 34609 33371 34667 33377
rect 34609 33337 34621 33371
rect 34655 33368 34667 33371
rect 37277 33371 37335 33377
rect 37277 33368 37289 33371
rect 34655 33340 37289 33368
rect 34655 33337 34667 33340
rect 34609 33331 34667 33337
rect 37277 33337 37289 33340
rect 37323 33337 37335 33371
rect 37277 33331 37335 33337
rect 26418 33300 26424 33312
rect 22888 33272 26004 33300
rect 26379 33272 26424 33300
rect 22888 33260 22894 33272
rect 26418 33260 26424 33272
rect 26476 33260 26482 33312
rect 26970 33260 26976 33312
rect 27028 33300 27034 33312
rect 29549 33303 29607 33309
rect 29549 33300 29561 33303
rect 27028 33272 29561 33300
rect 27028 33260 27034 33272
rect 29549 33269 29561 33272
rect 29595 33300 29607 33303
rect 29822 33300 29828 33312
rect 29595 33272 29828 33300
rect 29595 33269 29607 33272
rect 29549 33263 29607 33269
rect 29822 33260 29828 33272
rect 29880 33260 29886 33312
rect 36446 33300 36452 33312
rect 36407 33272 36452 33300
rect 36446 33260 36452 33272
rect 36504 33260 36510 33312
rect 37458 33300 37464 33312
rect 37419 33272 37464 33300
rect 37458 33260 37464 33272
rect 37516 33260 37522 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 15378 33096 15384 33108
rect 15339 33068 15384 33096
rect 15378 33056 15384 33068
rect 15436 33056 15442 33108
rect 16850 33056 16856 33108
rect 16908 33096 16914 33108
rect 17313 33099 17371 33105
rect 17313 33096 17325 33099
rect 16908 33068 17325 33096
rect 16908 33056 16914 33068
rect 17313 33065 17325 33068
rect 17359 33065 17371 33099
rect 17313 33059 17371 33065
rect 32398 33056 32404 33108
rect 32456 33096 32462 33108
rect 33045 33099 33103 33105
rect 33045 33096 33057 33099
rect 32456 33068 33057 33096
rect 32456 33056 32462 33068
rect 33045 33065 33057 33068
rect 33091 33096 33103 33099
rect 33134 33096 33140 33108
rect 33091 33068 33140 33096
rect 33091 33065 33103 33068
rect 33045 33059 33103 33065
rect 33134 33056 33140 33068
rect 33192 33056 33198 33108
rect 37550 33096 37556 33108
rect 37511 33068 37556 33096
rect 37550 33056 37556 33068
rect 37608 33056 37614 33108
rect 16868 32960 16896 33056
rect 18598 32960 18604 32972
rect 15580 32932 16896 32960
rect 17512 32932 18604 32960
rect 15580 32904 15608 32932
rect 15562 32892 15568 32904
rect 15475 32864 15568 32892
rect 15562 32852 15568 32864
rect 15620 32852 15626 32904
rect 15654 32852 15660 32904
rect 15712 32892 15718 32904
rect 17512 32901 17540 32932
rect 18598 32920 18604 32932
rect 18656 32920 18662 32972
rect 20990 32920 20996 32972
rect 21048 32960 21054 32972
rect 30193 32963 30251 32969
rect 30193 32960 30205 32963
rect 21048 32932 30205 32960
rect 21048 32920 21054 32932
rect 30193 32929 30205 32932
rect 30239 32960 30251 32963
rect 30239 32932 32260 32960
rect 30239 32929 30251 32932
rect 30193 32923 30251 32929
rect 32232 32904 32260 32932
rect 34514 32920 34520 32972
rect 34572 32960 34578 32972
rect 34701 32963 34759 32969
rect 34701 32960 34713 32963
rect 34572 32932 34713 32960
rect 34572 32920 34578 32932
rect 34701 32929 34713 32932
rect 34747 32929 34759 32963
rect 34701 32923 34759 32929
rect 34977 32963 35035 32969
rect 34977 32929 34989 32963
rect 35023 32960 35035 32963
rect 35802 32960 35808 32972
rect 35023 32932 35808 32960
rect 35023 32929 35035 32932
rect 34977 32923 35035 32929
rect 35802 32920 35808 32932
rect 35860 32920 35866 32972
rect 36170 32960 36176 32972
rect 36131 32932 36176 32960
rect 36170 32920 36176 32932
rect 36228 32920 36234 32972
rect 17497 32895 17555 32901
rect 15712 32864 15757 32892
rect 15712 32852 15718 32864
rect 17497 32861 17509 32895
rect 17543 32861 17555 32895
rect 17954 32892 17960 32904
rect 17915 32864 17960 32892
rect 17497 32855 17555 32861
rect 17954 32852 17960 32864
rect 18012 32852 18018 32904
rect 23658 32852 23664 32904
rect 23716 32892 23722 32904
rect 23753 32895 23811 32901
rect 23753 32892 23765 32895
rect 23716 32864 23765 32892
rect 23716 32852 23722 32864
rect 23753 32861 23765 32864
rect 23799 32861 23811 32895
rect 23753 32855 23811 32861
rect 30374 32852 30380 32904
rect 30432 32892 30438 32904
rect 30469 32895 30527 32901
rect 30469 32892 30481 32895
rect 30432 32864 30481 32892
rect 30432 32852 30438 32864
rect 30469 32861 30481 32864
rect 30515 32861 30527 32895
rect 30469 32855 30527 32861
rect 32033 32895 32091 32901
rect 32033 32861 32045 32895
rect 32079 32861 32091 32895
rect 32214 32892 32220 32904
rect 32175 32864 32220 32892
rect 32033 32855 32091 32861
rect 16942 32784 16948 32836
rect 17000 32824 17006 32836
rect 18141 32827 18199 32833
rect 18141 32824 18153 32827
rect 17000 32796 18153 32824
rect 17000 32784 17006 32796
rect 18141 32793 18153 32796
rect 18187 32793 18199 32827
rect 32048 32824 32076 32855
rect 32214 32852 32220 32864
rect 32272 32852 32278 32904
rect 36446 32901 36452 32904
rect 32401 32895 32459 32901
rect 32401 32861 32413 32895
rect 32447 32892 32459 32895
rect 32861 32895 32919 32901
rect 32861 32892 32873 32895
rect 32447 32864 32873 32892
rect 32447 32861 32459 32864
rect 32401 32855 32459 32861
rect 32861 32861 32873 32864
rect 32907 32861 32919 32895
rect 36440 32892 36452 32901
rect 36407 32864 36452 32892
rect 32861 32855 32919 32861
rect 36440 32855 36452 32864
rect 36446 32852 36452 32855
rect 36504 32852 36510 32904
rect 33226 32824 33232 32836
rect 32048 32796 33232 32824
rect 18141 32787 18199 32793
rect 33226 32784 33232 32796
rect 33284 32784 33290 32836
rect 18325 32759 18383 32765
rect 18325 32725 18337 32759
rect 18371 32756 18383 32759
rect 18506 32756 18512 32768
rect 18371 32728 18512 32756
rect 18371 32725 18383 32728
rect 18325 32719 18383 32725
rect 18506 32716 18512 32728
rect 18564 32716 18570 32768
rect 23658 32756 23664 32768
rect 23619 32728 23664 32756
rect 23658 32716 23664 32728
rect 23716 32716 23722 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 15654 32552 15660 32564
rect 15615 32524 15660 32552
rect 15654 32512 15660 32524
rect 15712 32552 15718 32564
rect 16666 32552 16672 32564
rect 15712 32524 16672 32552
rect 15712 32512 15718 32524
rect 16666 32512 16672 32524
rect 16724 32552 16730 32564
rect 16945 32555 17003 32561
rect 16945 32552 16957 32555
rect 16724 32524 16957 32552
rect 16724 32512 16730 32524
rect 16945 32521 16957 32524
rect 16991 32521 17003 32555
rect 16945 32515 17003 32521
rect 23477 32555 23535 32561
rect 23477 32521 23489 32555
rect 23523 32552 23535 32555
rect 23566 32552 23572 32564
rect 23523 32524 23572 32552
rect 23523 32521 23535 32524
rect 23477 32515 23535 32521
rect 23566 32512 23572 32524
rect 23624 32552 23630 32564
rect 24305 32555 24363 32561
rect 24305 32552 24317 32555
rect 23624 32524 24317 32552
rect 23624 32512 23630 32524
rect 24305 32521 24317 32524
rect 24351 32521 24363 32555
rect 24305 32515 24363 32521
rect 30653 32555 30711 32561
rect 30653 32521 30665 32555
rect 30699 32552 30711 32555
rect 30926 32552 30932 32564
rect 30699 32524 30932 32552
rect 30699 32521 30711 32524
rect 30653 32515 30711 32521
rect 30926 32512 30932 32524
rect 30984 32512 30990 32564
rect 37274 32552 37280 32564
rect 37235 32524 37280 32552
rect 37274 32512 37280 32524
rect 37332 32512 37338 32564
rect 15194 32484 15200 32496
rect 14292 32456 15200 32484
rect 14292 32425 14320 32456
rect 15194 32444 15200 32456
rect 15252 32484 15258 32496
rect 23014 32484 23020 32496
rect 15252 32456 18276 32484
rect 15252 32444 15258 32456
rect 14550 32425 14556 32428
rect 14277 32419 14335 32425
rect 14277 32385 14289 32419
rect 14323 32385 14335 32419
rect 14277 32379 14335 32385
rect 14544 32379 14556 32425
rect 14608 32416 14614 32428
rect 14608 32388 14644 32416
rect 14550 32376 14556 32379
rect 14608 32376 14614 32388
rect 16758 32376 16764 32428
rect 16816 32416 16822 32428
rect 16853 32419 16911 32425
rect 16853 32416 16865 32419
rect 16816 32388 16865 32416
rect 16816 32376 16822 32388
rect 16853 32385 16865 32388
rect 16899 32385 16911 32419
rect 17034 32416 17040 32428
rect 16995 32388 17040 32416
rect 16853 32379 16911 32385
rect 17034 32376 17040 32388
rect 17092 32376 17098 32428
rect 18248 32425 18276 32456
rect 22112 32456 23020 32484
rect 18233 32419 18291 32425
rect 18233 32385 18245 32419
rect 18279 32385 18291 32419
rect 18233 32379 18291 32385
rect 18322 32376 18328 32428
rect 18380 32416 18386 32428
rect 18489 32419 18547 32425
rect 18489 32416 18501 32419
rect 18380 32388 18501 32416
rect 18380 32376 18386 32388
rect 18489 32385 18501 32388
rect 18535 32385 18547 32419
rect 18489 32379 18547 32385
rect 20441 32419 20499 32425
rect 20441 32385 20453 32419
rect 20487 32416 20499 32419
rect 20990 32416 20996 32428
rect 20487 32388 20996 32416
rect 20487 32385 20499 32388
rect 20441 32379 20499 32385
rect 20990 32376 20996 32388
rect 21048 32376 21054 32428
rect 22112 32425 22140 32456
rect 23014 32444 23020 32456
rect 23072 32444 23078 32496
rect 27522 32444 27528 32496
rect 27580 32484 27586 32496
rect 28169 32487 28227 32493
rect 28169 32484 28181 32487
rect 27580 32456 28181 32484
rect 27580 32444 27586 32456
rect 28169 32453 28181 32456
rect 28215 32453 28227 32487
rect 28169 32447 28227 32453
rect 30285 32487 30343 32493
rect 30285 32453 30297 32487
rect 30331 32484 30343 32487
rect 30374 32484 30380 32496
rect 30331 32456 30380 32484
rect 30331 32453 30343 32456
rect 30285 32447 30343 32453
rect 30374 32444 30380 32456
rect 30432 32444 30438 32496
rect 30466 32444 30472 32496
rect 30524 32493 30530 32496
rect 30524 32487 30543 32493
rect 30531 32453 30543 32487
rect 31294 32484 31300 32496
rect 31255 32456 31300 32484
rect 30524 32447 30543 32453
rect 30524 32444 30530 32447
rect 31294 32444 31300 32456
rect 31352 32444 31358 32496
rect 32214 32444 32220 32496
rect 32272 32484 32278 32496
rect 32309 32487 32367 32493
rect 32309 32484 32321 32487
rect 32272 32456 32321 32484
rect 32272 32444 32278 32456
rect 32309 32453 32321 32456
rect 32355 32453 32367 32487
rect 32309 32447 32367 32453
rect 33312 32487 33370 32493
rect 33312 32453 33324 32487
rect 33358 32484 33370 32487
rect 33502 32484 33508 32496
rect 33358 32456 33508 32484
rect 33358 32453 33370 32456
rect 33312 32447 33370 32453
rect 33502 32444 33508 32456
rect 33560 32444 33566 32496
rect 35802 32444 35808 32496
rect 35860 32484 35866 32496
rect 35860 32456 37504 32484
rect 35860 32444 35866 32456
rect 22097 32419 22155 32425
rect 22097 32385 22109 32419
rect 22143 32385 22155 32419
rect 22097 32379 22155 32385
rect 22364 32419 22422 32425
rect 22364 32385 22376 32419
rect 22410 32416 22422 32419
rect 23198 32416 23204 32428
rect 22410 32388 23204 32416
rect 22410 32385 22422 32388
rect 22364 32379 22422 32385
rect 23198 32376 23204 32388
rect 23256 32376 23262 32428
rect 24121 32419 24179 32425
rect 24121 32385 24133 32419
rect 24167 32385 24179 32419
rect 24121 32379 24179 32385
rect 24397 32419 24455 32425
rect 24397 32385 24409 32419
rect 24443 32416 24455 32419
rect 24854 32416 24860 32428
rect 24443 32388 24860 32416
rect 24443 32385 24455 32388
rect 24397 32379 24455 32385
rect 20622 32348 20628 32360
rect 19628 32320 20628 32348
rect 16574 32240 16580 32292
rect 16632 32280 16638 32292
rect 19628 32289 19656 32320
rect 20622 32308 20628 32320
rect 20680 32308 20686 32360
rect 16669 32283 16727 32289
rect 16669 32280 16681 32283
rect 16632 32252 16681 32280
rect 16632 32240 16638 32252
rect 16669 32249 16681 32252
rect 16715 32249 16727 32283
rect 16669 32243 16727 32249
rect 19613 32283 19671 32289
rect 19613 32249 19625 32283
rect 19659 32249 19671 32283
rect 24136 32280 24164 32379
rect 24854 32376 24860 32388
rect 24912 32376 24918 32428
rect 25317 32419 25375 32425
rect 25317 32385 25329 32419
rect 25363 32385 25375 32419
rect 25317 32379 25375 32385
rect 25332 32348 25360 32379
rect 25406 32376 25412 32428
rect 25464 32416 25470 32428
rect 25593 32419 25651 32425
rect 25464 32388 25509 32416
rect 25464 32376 25470 32388
rect 25593 32385 25605 32419
rect 25639 32416 25651 32419
rect 25866 32416 25872 32428
rect 25639 32388 25872 32416
rect 25639 32385 25651 32388
rect 25593 32379 25651 32385
rect 25866 32376 25872 32388
rect 25924 32376 25930 32428
rect 27985 32419 28043 32425
rect 27985 32385 27997 32419
rect 28031 32385 28043 32419
rect 27985 32379 28043 32385
rect 28261 32419 28319 32425
rect 28261 32385 28273 32419
rect 28307 32385 28319 32419
rect 28261 32379 28319 32385
rect 28353 32419 28411 32425
rect 28353 32385 28365 32419
rect 28399 32416 28411 32419
rect 28902 32416 28908 32428
rect 28399 32388 28908 32416
rect 28399 32385 28411 32388
rect 28353 32379 28411 32385
rect 25774 32348 25780 32360
rect 25332 32320 25780 32348
rect 25774 32308 25780 32320
rect 25832 32308 25838 32360
rect 27890 32280 27896 32292
rect 24136 32252 27896 32280
rect 19613 32243 19671 32249
rect 27890 32240 27896 32252
rect 27948 32240 27954 32292
rect 28000 32280 28028 32379
rect 28276 32348 28304 32379
rect 28902 32376 28908 32388
rect 28960 32376 28966 32428
rect 31481 32419 31539 32425
rect 31481 32385 31493 32419
rect 31527 32416 31539 32419
rect 32490 32416 32496 32428
rect 31527 32388 32496 32416
rect 31527 32385 31539 32388
rect 31481 32379 31539 32385
rect 32490 32376 32496 32388
rect 32548 32376 32554 32428
rect 36096 32425 36124 32456
rect 35253 32419 35311 32425
rect 35253 32385 35265 32419
rect 35299 32416 35311 32419
rect 35897 32419 35955 32425
rect 35897 32416 35909 32419
rect 35299 32388 35909 32416
rect 35299 32385 35311 32388
rect 35253 32379 35311 32385
rect 35897 32385 35909 32388
rect 35943 32385 35955 32419
rect 35897 32379 35955 32385
rect 36081 32419 36139 32425
rect 36081 32385 36093 32419
rect 36127 32385 36139 32419
rect 36262 32416 36268 32428
rect 36223 32388 36268 32416
rect 36081 32379 36139 32385
rect 36262 32376 36268 32388
rect 36320 32376 36326 32428
rect 37476 32425 37504 32456
rect 37461 32419 37519 32425
rect 37461 32385 37473 32419
rect 37507 32385 37519 32419
rect 37461 32379 37519 32385
rect 37645 32419 37703 32425
rect 37645 32385 37657 32419
rect 37691 32416 37703 32419
rect 37734 32416 37740 32428
rect 37691 32388 37740 32416
rect 37691 32385 37703 32388
rect 37645 32379 37703 32385
rect 37734 32376 37740 32388
rect 37792 32376 37798 32428
rect 28442 32348 28448 32360
rect 28276 32320 28448 32348
rect 28442 32308 28448 32320
rect 28500 32348 28506 32360
rect 29822 32348 29828 32360
rect 28500 32320 29828 32348
rect 28500 32308 28506 32320
rect 29822 32308 29828 32320
rect 29880 32308 29886 32360
rect 32030 32308 32036 32360
rect 32088 32348 32094 32360
rect 33045 32351 33103 32357
rect 33045 32348 33057 32351
rect 32088 32320 33057 32348
rect 32088 32308 32094 32320
rect 33045 32317 33057 32320
rect 33091 32317 33103 32351
rect 33045 32311 33103 32317
rect 28258 32280 28264 32292
rect 28000 32252 28264 32280
rect 28258 32240 28264 32252
rect 28316 32280 28322 32292
rect 28626 32280 28632 32292
rect 28316 32252 28632 32280
rect 28316 32240 28322 32252
rect 28626 32240 28632 32252
rect 28684 32240 28690 32292
rect 17221 32215 17279 32221
rect 17221 32181 17233 32215
rect 17267 32212 17279 32215
rect 18230 32212 18236 32224
rect 17267 32184 18236 32212
rect 17267 32181 17279 32184
rect 17221 32175 17279 32181
rect 18230 32172 18236 32184
rect 18288 32172 18294 32224
rect 20254 32212 20260 32224
rect 20215 32184 20260 32212
rect 20254 32172 20260 32184
rect 20312 32172 20318 32224
rect 23934 32212 23940 32224
rect 23895 32184 23940 32212
rect 23934 32172 23940 32184
rect 23992 32172 23998 32224
rect 25777 32215 25835 32221
rect 25777 32181 25789 32215
rect 25823 32212 25835 32215
rect 27154 32212 27160 32224
rect 25823 32184 27160 32212
rect 25823 32181 25835 32184
rect 25777 32175 25835 32181
rect 27154 32172 27160 32184
rect 27212 32172 27218 32224
rect 28350 32172 28356 32224
rect 28408 32212 28414 32224
rect 28537 32215 28595 32221
rect 28537 32212 28549 32215
rect 28408 32184 28549 32212
rect 28408 32172 28414 32184
rect 28537 32181 28549 32184
rect 28583 32181 28595 32215
rect 28537 32175 28595 32181
rect 30374 32172 30380 32224
rect 30432 32212 30438 32224
rect 30469 32215 30527 32221
rect 30469 32212 30481 32215
rect 30432 32184 30481 32212
rect 30432 32172 30438 32184
rect 30469 32181 30481 32184
rect 30515 32181 30527 32215
rect 30469 32175 30527 32181
rect 33226 32172 33232 32224
rect 33284 32212 33290 32224
rect 34425 32215 34483 32221
rect 34425 32212 34437 32215
rect 33284 32184 34437 32212
rect 33284 32172 33290 32184
rect 34425 32181 34437 32184
rect 34471 32181 34483 32215
rect 35434 32212 35440 32224
rect 35395 32184 35440 32212
rect 34425 32175 34483 32181
rect 35434 32172 35440 32184
rect 35492 32172 35498 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 14550 31968 14556 32020
rect 14608 32008 14614 32020
rect 14737 32011 14795 32017
rect 14737 32008 14749 32011
rect 14608 31980 14749 32008
rect 14608 31968 14614 31980
rect 14737 31977 14749 31980
rect 14783 31977 14795 32011
rect 16758 32008 16764 32020
rect 16719 31980 16764 32008
rect 14737 31971 14795 31977
rect 16758 31968 16764 31980
rect 16816 31968 16822 32020
rect 16942 32008 16948 32020
rect 16903 31980 16948 32008
rect 16942 31968 16948 31980
rect 17000 31968 17006 32020
rect 18049 32011 18107 32017
rect 18049 31977 18061 32011
rect 18095 32008 18107 32011
rect 18322 32008 18328 32020
rect 18095 31980 18328 32008
rect 18095 31977 18107 31980
rect 18049 31971 18107 31977
rect 18322 31968 18328 31980
rect 18380 31968 18386 32020
rect 18598 31968 18604 32020
rect 18656 32008 18662 32020
rect 22002 32008 22008 32020
rect 18656 31980 22008 32008
rect 18656 31968 18662 31980
rect 22002 31968 22008 31980
rect 22060 31968 22066 32020
rect 23198 32008 23204 32020
rect 23159 31980 23204 32008
rect 23198 31968 23204 31980
rect 23256 31968 23262 32020
rect 26053 32011 26111 32017
rect 26053 31977 26065 32011
rect 26099 32008 26111 32011
rect 26234 32008 26240 32020
rect 26099 31980 26240 32008
rect 26099 31977 26111 31980
rect 26053 31971 26111 31977
rect 26234 31968 26240 31980
rect 26292 32008 26298 32020
rect 30742 32008 30748 32020
rect 26292 31980 30748 32008
rect 26292 31968 26298 31980
rect 30742 31968 30748 31980
rect 30800 31968 30806 32020
rect 30926 32008 30932 32020
rect 30887 31980 30932 32008
rect 30926 31968 30932 31980
rect 30984 31968 30990 32020
rect 33965 32011 34023 32017
rect 31726 31980 33272 32008
rect 17034 31940 17040 31952
rect 15764 31912 17040 31940
rect 14921 31807 14979 31813
rect 14921 31773 14933 31807
rect 14967 31804 14979 31807
rect 15381 31807 15439 31813
rect 15381 31804 15393 31807
rect 14967 31776 15393 31804
rect 14967 31773 14979 31776
rect 14921 31767 14979 31773
rect 15381 31773 15393 31776
rect 15427 31773 15439 31807
rect 15562 31804 15568 31816
rect 15523 31776 15568 31804
rect 15381 31767 15439 31773
rect 15562 31764 15568 31776
rect 15620 31764 15626 31816
rect 15764 31813 15792 31912
rect 16500 31813 16528 31912
rect 17034 31900 17040 31912
rect 17092 31900 17098 31952
rect 19337 31943 19395 31949
rect 19337 31940 19349 31943
rect 18708 31912 19349 31940
rect 18708 31884 18736 31912
rect 19337 31909 19349 31912
rect 19383 31909 19395 31943
rect 20714 31940 20720 31952
rect 19337 31903 19395 31909
rect 19444 31912 20720 31940
rect 16666 31872 16672 31884
rect 16627 31844 16672 31872
rect 16666 31832 16672 31844
rect 16724 31832 16730 31884
rect 18414 31872 18420 31884
rect 18340 31844 18420 31872
rect 15749 31807 15807 31813
rect 15749 31773 15761 31807
rect 15795 31773 15807 31807
rect 15749 31767 15807 31773
rect 16485 31807 16543 31813
rect 16485 31773 16497 31807
rect 16531 31773 16543 31807
rect 16485 31767 16543 31773
rect 16761 31807 16819 31813
rect 16761 31773 16773 31807
rect 16807 31773 16819 31807
rect 18230 31804 18236 31816
rect 18191 31776 18236 31804
rect 16761 31767 16819 31773
rect 16666 31696 16672 31748
rect 16724 31736 16730 31748
rect 16776 31736 16804 31767
rect 18230 31764 18236 31776
rect 18288 31764 18294 31816
rect 18340 31813 18368 31844
rect 18414 31832 18420 31844
rect 18472 31832 18478 31884
rect 18690 31872 18696 31884
rect 18603 31844 18696 31872
rect 18690 31832 18696 31844
rect 18748 31832 18754 31884
rect 18325 31807 18383 31813
rect 18325 31773 18337 31807
rect 18371 31773 18383 31807
rect 18325 31767 18383 31773
rect 18506 31764 18512 31816
rect 18564 31813 18570 31816
rect 18564 31807 18593 31813
rect 18581 31773 18593 31807
rect 19444 31804 19472 31912
rect 20714 31900 20720 31912
rect 20772 31900 20778 31952
rect 20901 31943 20959 31949
rect 20901 31909 20913 31943
rect 20947 31940 20959 31943
rect 21266 31940 21272 31952
rect 20947 31912 21272 31940
rect 20947 31909 20959 31912
rect 20901 31903 20959 31909
rect 21266 31900 21272 31912
rect 21324 31900 21330 31952
rect 22738 31900 22744 31952
rect 22796 31940 22802 31952
rect 23014 31940 23020 31952
rect 22796 31912 23020 31940
rect 22796 31900 22802 31912
rect 23014 31900 23020 31912
rect 23072 31900 23078 31952
rect 27338 31900 27344 31952
rect 27396 31940 27402 31952
rect 31726 31940 31754 31980
rect 27396 31912 31754 31940
rect 32033 31943 32091 31949
rect 27396 31900 27402 31912
rect 32033 31909 32045 31943
rect 32079 31940 32091 31943
rect 32490 31940 32496 31952
rect 32079 31912 32496 31940
rect 32079 31909 32091 31912
rect 32033 31903 32091 31909
rect 32490 31900 32496 31912
rect 32548 31940 32554 31952
rect 33244 31940 33272 31980
rect 33965 31977 33977 32011
rect 34011 32008 34023 32011
rect 34422 32008 34428 32020
rect 34011 31980 34428 32008
rect 34011 31977 34023 31980
rect 33965 31971 34023 31977
rect 34422 31968 34428 31980
rect 34480 31968 34486 32020
rect 35342 31940 35348 31952
rect 32548 31912 33180 31940
rect 33244 31912 35348 31940
rect 32548 31900 32554 31912
rect 20622 31872 20628 31884
rect 20583 31844 20628 31872
rect 20622 31832 20628 31844
rect 20680 31832 20686 31884
rect 20990 31832 20996 31884
rect 21048 31872 21054 31884
rect 21085 31875 21143 31881
rect 21085 31872 21097 31875
rect 21048 31844 21097 31872
rect 21048 31832 21054 31844
rect 21085 31841 21097 31844
rect 21131 31841 21143 31875
rect 23382 31872 23388 31884
rect 21085 31835 21143 31841
rect 22940 31844 23388 31872
rect 18564 31767 18593 31773
rect 18708 31776 19472 31804
rect 19521 31807 19579 31813
rect 18564 31764 18570 31767
rect 16724 31708 16804 31736
rect 18417 31739 18475 31745
rect 16724 31696 16730 31708
rect 18417 31705 18429 31739
rect 18463 31736 18475 31739
rect 18708 31736 18736 31776
rect 19521 31773 19533 31807
rect 19567 31804 19579 31807
rect 20254 31804 20260 31816
rect 19567 31776 20260 31804
rect 19567 31773 19579 31776
rect 19521 31767 19579 31773
rect 20254 31764 20260 31776
rect 20312 31764 20318 31816
rect 22940 31813 22968 31844
rect 23382 31832 23388 31844
rect 23440 31832 23446 31884
rect 24857 31875 24915 31881
rect 24857 31841 24869 31875
rect 24903 31872 24915 31875
rect 30374 31872 30380 31884
rect 24903 31844 30380 31872
rect 24903 31841 24915 31844
rect 24857 31835 24915 31841
rect 30374 31832 30380 31844
rect 30432 31872 30438 31884
rect 30745 31875 30803 31881
rect 30745 31872 30757 31875
rect 30432 31844 30757 31872
rect 30432 31832 30438 31844
rect 30745 31841 30757 31844
rect 30791 31841 30803 31875
rect 30745 31835 30803 31841
rect 22925 31807 22983 31813
rect 22925 31773 22937 31807
rect 22971 31773 22983 31807
rect 22925 31767 22983 31773
rect 23017 31807 23075 31813
rect 23017 31773 23029 31807
rect 23063 31804 23075 31807
rect 23201 31807 23259 31813
rect 23063 31776 23152 31804
rect 23063 31773 23075 31776
rect 23017 31767 23075 31773
rect 18463 31708 18736 31736
rect 23124 31736 23152 31776
rect 23201 31773 23213 31807
rect 23247 31804 23259 31807
rect 23934 31804 23940 31816
rect 23247 31776 23940 31804
rect 23247 31773 23259 31776
rect 23201 31767 23259 31773
rect 23934 31764 23940 31776
rect 23992 31764 23998 31816
rect 24578 31804 24584 31816
rect 24044 31776 24584 31804
rect 23658 31736 23664 31748
rect 23124 31708 23664 31736
rect 18463 31705 18475 31708
rect 18417 31699 18475 31705
rect 23658 31696 23664 31708
rect 23716 31736 23722 31748
rect 24044 31736 24072 31776
rect 24578 31764 24584 31776
rect 24636 31764 24642 31816
rect 24673 31807 24731 31813
rect 24673 31773 24685 31807
rect 24719 31804 24731 31807
rect 25038 31804 25044 31816
rect 24719 31776 25044 31804
rect 24719 31773 24731 31776
rect 24673 31767 24731 31773
rect 25038 31764 25044 31776
rect 25096 31764 25102 31816
rect 27338 31804 27344 31816
rect 27299 31776 27344 31804
rect 27338 31764 27344 31776
rect 27396 31764 27402 31816
rect 28902 31764 28908 31816
rect 28960 31804 28966 31816
rect 29546 31804 29552 31816
rect 28960 31776 29408 31804
rect 29507 31776 29552 31804
rect 28960 31764 28966 31776
rect 23716 31708 24072 31736
rect 29380 31736 29408 31776
rect 29546 31764 29552 31776
rect 29604 31764 29610 31816
rect 29733 31807 29791 31813
rect 29733 31804 29745 31807
rect 29656 31776 29745 31804
rect 29656 31736 29684 31776
rect 29733 31773 29745 31776
rect 29779 31773 29791 31807
rect 29825 31807 29883 31813
rect 29825 31794 29837 31807
rect 29871 31794 29883 31807
rect 29733 31767 29791 31773
rect 29822 31742 29828 31794
rect 29880 31742 29886 31794
rect 29914 31764 29920 31816
rect 29972 31804 29978 31816
rect 30101 31807 30159 31813
rect 29972 31776 30017 31804
rect 29972 31764 29978 31776
rect 30101 31773 30113 31807
rect 30147 31804 30159 31807
rect 30190 31804 30196 31816
rect 30147 31776 30196 31804
rect 30147 31773 30159 31776
rect 30101 31767 30159 31773
rect 30190 31764 30196 31776
rect 30248 31764 30254 31816
rect 31205 31807 31263 31813
rect 31205 31773 31217 31807
rect 31251 31804 31263 31807
rect 31294 31804 31300 31816
rect 31251 31776 31300 31804
rect 31251 31773 31263 31776
rect 31205 31767 31263 31773
rect 31294 31764 31300 31776
rect 31352 31764 31358 31816
rect 31754 31764 31760 31816
rect 31812 31804 31818 31816
rect 33152 31813 33180 31912
rect 35342 31900 35348 31912
rect 35400 31900 35406 31952
rect 36449 31875 36507 31881
rect 36449 31841 36461 31875
rect 36495 31872 36507 31875
rect 37458 31872 37464 31884
rect 36495 31844 37464 31872
rect 36495 31841 36507 31844
rect 36449 31835 36507 31841
rect 37458 31832 37464 31844
rect 37516 31832 37522 31884
rect 38102 31872 38108 31884
rect 38063 31844 38108 31872
rect 38102 31832 38108 31844
rect 38160 31832 38166 31884
rect 32125 31807 32183 31813
rect 32125 31804 32137 31807
rect 31812 31776 32137 31804
rect 31812 31764 31818 31776
rect 32125 31773 32137 31776
rect 32171 31773 32183 31807
rect 33045 31807 33103 31813
rect 33045 31780 33057 31807
rect 32125 31767 32183 31773
rect 32968 31773 33057 31780
rect 33091 31773 33103 31807
rect 32968 31767 33103 31773
rect 33137 31807 33195 31813
rect 33137 31773 33149 31807
rect 33183 31773 33195 31807
rect 33137 31767 33195 31773
rect 32968 31752 33088 31767
rect 33226 31764 33232 31816
rect 33284 31764 33290 31816
rect 33321 31807 33379 31813
rect 33321 31773 33333 31807
rect 33367 31804 33379 31807
rect 33781 31807 33839 31813
rect 33781 31804 33793 31807
rect 33367 31776 33793 31804
rect 33367 31773 33379 31776
rect 33321 31767 33379 31773
rect 33781 31773 33793 31776
rect 33827 31773 33839 31807
rect 33781 31767 33839 31773
rect 35805 31807 35863 31813
rect 35805 31773 35817 31807
rect 35851 31804 35863 31807
rect 36265 31807 36323 31813
rect 36265 31804 36277 31807
rect 35851 31776 36277 31804
rect 35851 31773 35863 31776
rect 35805 31767 35863 31773
rect 36265 31773 36277 31776
rect 36311 31773 36323 31807
rect 36265 31767 36323 31773
rect 29380 31708 29684 31736
rect 23716 31696 23722 31708
rect 24857 31671 24915 31677
rect 24857 31637 24869 31671
rect 24903 31668 24915 31671
rect 26050 31668 26056 31680
rect 24903 31640 26056 31668
rect 24903 31637 24915 31640
rect 24857 31631 24915 31637
rect 26050 31628 26056 31640
rect 26108 31628 26114 31680
rect 29454 31628 29460 31680
rect 29512 31668 29518 31680
rect 30285 31671 30343 31677
rect 30285 31668 30297 31671
rect 29512 31640 30297 31668
rect 29512 31628 29518 31640
rect 30285 31637 30297 31640
rect 30331 31637 30343 31671
rect 32968 31668 32996 31752
rect 33244 31668 33272 31764
rect 32968 31640 33272 31668
rect 30285 31631 30343 31637
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 10962 31424 10968 31476
rect 11020 31464 11026 31476
rect 11020 31436 25084 31464
rect 11020 31424 11026 31436
rect 18690 31405 18696 31408
rect 18684 31396 18696 31405
rect 15672 31368 16896 31396
rect 18651 31368 18696 31396
rect 15562 31328 15568 31340
rect 15523 31300 15568 31328
rect 15562 31288 15568 31300
rect 15620 31328 15626 31340
rect 15672 31328 15700 31368
rect 15620 31300 15700 31328
rect 15749 31331 15807 31337
rect 15620 31288 15626 31300
rect 15749 31297 15761 31331
rect 15795 31328 15807 31331
rect 16758 31328 16764 31340
rect 15795 31300 16764 31328
rect 15795 31297 15807 31300
rect 15749 31291 15807 31297
rect 16758 31288 16764 31300
rect 16816 31288 16822 31340
rect 16868 31337 16896 31368
rect 18684 31359 18696 31368
rect 18690 31356 18696 31359
rect 18748 31356 18754 31408
rect 20070 31356 20076 31408
rect 20128 31396 20134 31408
rect 20901 31399 20959 31405
rect 20901 31396 20913 31399
rect 20128 31368 20913 31396
rect 20128 31356 20134 31368
rect 20901 31365 20913 31368
rect 20947 31365 20959 31399
rect 20901 31359 20959 31365
rect 21018 31399 21076 31405
rect 21018 31365 21030 31399
rect 21064 31396 21076 31399
rect 21266 31396 21272 31408
rect 21064 31368 21272 31396
rect 21064 31365 21076 31368
rect 21018 31359 21076 31365
rect 16853 31331 16911 31337
rect 16853 31297 16865 31331
rect 16899 31297 16911 31331
rect 16853 31291 16911 31297
rect 17037 31331 17095 31337
rect 17037 31297 17049 31331
rect 17083 31328 17095 31331
rect 17497 31331 17555 31337
rect 17497 31328 17509 31331
rect 17083 31300 17509 31328
rect 17083 31297 17095 31300
rect 17037 31291 17095 31297
rect 17497 31297 17509 31300
rect 17543 31297 17555 31331
rect 17497 31291 17555 31297
rect 20533 31331 20591 31337
rect 20533 31297 20545 31331
rect 20579 31328 20591 31331
rect 20622 31328 20628 31340
rect 20579 31300 20628 31328
rect 20579 31297 20591 31300
rect 20533 31291 20591 31297
rect 20622 31288 20628 31300
rect 20680 31288 20686 31340
rect 20916 31328 20944 31359
rect 21266 31356 21272 31368
rect 21324 31356 21330 31408
rect 23014 31405 23020 31408
rect 23008 31396 23020 31405
rect 22975 31368 23020 31396
rect 23008 31359 23020 31368
rect 23014 31356 23020 31359
rect 23072 31356 23078 31408
rect 21818 31328 21824 31340
rect 20916 31300 21824 31328
rect 21818 31288 21824 31300
rect 21876 31288 21882 31340
rect 24762 31328 24768 31340
rect 24136 31300 24768 31328
rect 16666 31260 16672 31272
rect 16627 31232 16672 31260
rect 16666 31220 16672 31232
rect 16724 31220 16730 31272
rect 18414 31260 18420 31272
rect 18375 31232 18420 31260
rect 18414 31220 18420 31232
rect 18472 31220 18478 31272
rect 20806 31260 20812 31272
rect 19812 31232 20812 31260
rect 19812 31201 19840 31232
rect 20806 31220 20812 31232
rect 20864 31220 20870 31272
rect 22462 31220 22468 31272
rect 22520 31260 22526 31272
rect 22741 31263 22799 31269
rect 22741 31260 22753 31263
rect 22520 31232 22753 31260
rect 22520 31220 22526 31232
rect 22741 31229 22753 31232
rect 22787 31229 22799 31263
rect 22741 31223 22799 31229
rect 24136 31201 24164 31300
rect 24762 31288 24768 31300
rect 24820 31328 24826 31340
rect 24857 31331 24915 31337
rect 24857 31328 24869 31331
rect 24820 31300 24869 31328
rect 24820 31288 24826 31300
rect 24857 31297 24869 31300
rect 24903 31297 24915 31331
rect 24857 31291 24915 31297
rect 25056 31260 25084 31436
rect 25222 31424 25228 31476
rect 25280 31424 25286 31476
rect 25406 31464 25412 31476
rect 25367 31436 25412 31464
rect 25406 31424 25412 31436
rect 25464 31424 25470 31476
rect 25774 31424 25780 31476
rect 25832 31464 25838 31476
rect 25869 31467 25927 31473
rect 25869 31464 25881 31467
rect 25832 31436 25881 31464
rect 25832 31424 25838 31436
rect 25869 31433 25881 31436
rect 25915 31433 25927 31467
rect 25869 31427 25927 31433
rect 26050 31424 26056 31476
rect 26108 31464 26114 31476
rect 26108 31436 26464 31464
rect 26108 31424 26114 31436
rect 25240 31396 25268 31424
rect 26145 31399 26203 31405
rect 26145 31396 26157 31399
rect 25148 31368 26157 31396
rect 25148 31337 25176 31368
rect 26145 31365 26157 31368
rect 26191 31365 26203 31399
rect 26145 31359 26203 31365
rect 25133 31331 25191 31337
rect 25133 31297 25145 31331
rect 25179 31297 25191 31331
rect 25133 31291 25191 31297
rect 25225 31331 25283 31337
rect 25225 31297 25237 31331
rect 25271 31328 25283 31331
rect 26050 31328 26056 31340
rect 25271 31300 26056 31328
rect 25271 31297 25283 31300
rect 25225 31291 25283 31297
rect 26050 31288 26056 31300
rect 26108 31288 26114 31340
rect 26237 31331 26295 31337
rect 26237 31297 26249 31331
rect 26283 31328 26295 31331
rect 26326 31328 26332 31340
rect 26283 31300 26332 31328
rect 26283 31297 26295 31300
rect 26237 31291 26295 31297
rect 26326 31288 26332 31300
rect 26384 31288 26390 31340
rect 26436 31337 26464 31436
rect 29270 31424 29276 31476
rect 29328 31464 29334 31476
rect 30006 31464 30012 31476
rect 29328 31436 30012 31464
rect 29328 31424 29334 31436
rect 28534 31356 28540 31408
rect 28592 31405 28598 31408
rect 28592 31396 28604 31405
rect 28592 31368 28637 31396
rect 28592 31359 28604 31368
rect 28592 31356 28598 31359
rect 26421 31331 26479 31337
rect 26421 31297 26433 31331
rect 26467 31297 26479 31331
rect 26421 31291 26479 31297
rect 27154 31288 27160 31340
rect 27212 31328 27218 31340
rect 28074 31328 28080 31340
rect 27212 31300 28080 31328
rect 27212 31288 27218 31300
rect 28074 31288 28080 31300
rect 28132 31288 28138 31340
rect 29454 31328 29460 31340
rect 29415 31300 29460 31328
rect 29454 31288 29460 31300
rect 29512 31288 29518 31340
rect 29564 31337 29592 31436
rect 30006 31424 30012 31436
rect 30064 31424 30070 31476
rect 30101 31467 30159 31473
rect 30101 31433 30113 31467
rect 30147 31464 30159 31467
rect 30374 31464 30380 31476
rect 30147 31436 30380 31464
rect 30147 31433 30159 31436
rect 30101 31427 30159 31433
rect 30374 31424 30380 31436
rect 30432 31424 30438 31476
rect 30926 31464 30932 31476
rect 30484 31436 30932 31464
rect 29825 31399 29883 31405
rect 29825 31365 29837 31399
rect 29871 31396 29883 31399
rect 30484 31396 30512 31436
rect 30926 31424 30932 31436
rect 30984 31424 30990 31476
rect 37458 31424 37464 31476
rect 37516 31464 37522 31476
rect 37553 31467 37611 31473
rect 37553 31464 37565 31467
rect 37516 31436 37565 31464
rect 37516 31424 37522 31436
rect 37553 31433 37565 31436
rect 37599 31433 37611 31467
rect 37553 31427 37611 31433
rect 29871 31368 30512 31396
rect 32140 31368 34100 31396
rect 29871 31365 29883 31368
rect 29825 31359 29883 31365
rect 29550 31331 29608 31337
rect 29550 31297 29562 31331
rect 29596 31297 29608 31331
rect 29550 31291 29608 31297
rect 29730 31288 29736 31340
rect 29788 31328 29794 31340
rect 29963 31331 30021 31337
rect 29788 31300 29833 31328
rect 29788 31288 29794 31300
rect 29963 31297 29975 31331
rect 30009 31328 30021 31331
rect 30653 31331 30711 31337
rect 30653 31328 30665 31331
rect 30009 31300 30665 31328
rect 30009 31297 30021 31300
rect 29963 31291 30021 31297
rect 30653 31297 30665 31300
rect 30699 31297 30711 31331
rect 30653 31291 30711 31297
rect 30745 31331 30803 31337
rect 30745 31297 30757 31331
rect 30791 31328 30803 31331
rect 31294 31328 31300 31340
rect 30791 31300 31300 31328
rect 30791 31297 30803 31300
rect 30745 31291 30803 31297
rect 31294 31288 31300 31300
rect 31352 31288 31358 31340
rect 31662 31288 31668 31340
rect 31720 31328 31726 31340
rect 32140 31337 32168 31368
rect 32398 31337 32404 31340
rect 32125 31331 32183 31337
rect 32125 31328 32137 31331
rect 31720 31300 32137 31328
rect 31720 31288 31726 31300
rect 32125 31297 32137 31300
rect 32171 31297 32183 31331
rect 32392 31328 32404 31337
rect 32359 31300 32404 31328
rect 32125 31291 32183 31297
rect 32392 31291 32404 31300
rect 32398 31288 32404 31291
rect 32456 31288 32462 31340
rect 34072 31272 34100 31368
rect 35434 31356 35440 31408
rect 35492 31396 35498 31408
rect 35590 31399 35648 31405
rect 35590 31396 35602 31399
rect 35492 31368 35602 31396
rect 35492 31356 35498 31368
rect 35590 31365 35602 31368
rect 35636 31365 35648 31399
rect 35590 31359 35648 31365
rect 37461 31331 37519 31337
rect 37461 31297 37473 31331
rect 37507 31328 37519 31331
rect 37550 31328 37556 31340
rect 37507 31300 37556 31328
rect 37507 31297 37519 31300
rect 37461 31291 37519 31297
rect 37550 31288 37556 31300
rect 37608 31288 37614 31340
rect 28813 31263 28871 31269
rect 25056 31232 27568 31260
rect 19797 31195 19855 31201
rect 19797 31161 19809 31195
rect 19843 31161 19855 31195
rect 19797 31155 19855 31161
rect 24121 31195 24179 31201
rect 24121 31161 24133 31195
rect 24167 31161 24179 31195
rect 24121 31155 24179 31161
rect 14274 31084 14280 31136
rect 14332 31124 14338 31136
rect 15381 31127 15439 31133
rect 15381 31124 15393 31127
rect 14332 31096 15393 31124
rect 14332 31084 14338 31096
rect 15381 31093 15393 31096
rect 15427 31093 15439 31127
rect 17678 31124 17684 31136
rect 17639 31096 17684 31124
rect 15381 31087 15439 31093
rect 17678 31084 17684 31096
rect 17736 31084 17742 31136
rect 21174 31124 21180 31136
rect 21135 31096 21180 31124
rect 21174 31084 21180 31096
rect 21232 31084 21238 31136
rect 24949 31127 25007 31133
rect 24949 31093 24961 31127
rect 24995 31124 25007 31127
rect 25498 31124 25504 31136
rect 24995 31096 25504 31124
rect 24995 31093 25007 31096
rect 24949 31087 25007 31093
rect 25498 31084 25504 31096
rect 25556 31084 25562 31136
rect 27430 31124 27436 31136
rect 27391 31096 27436 31124
rect 27430 31084 27436 31096
rect 27488 31084 27494 31136
rect 27540 31124 27568 31232
rect 28813 31229 28825 31263
rect 28859 31260 28871 31263
rect 32030 31260 32036 31272
rect 28859 31232 32036 31260
rect 28859 31229 28871 31232
rect 28813 31223 28871 31229
rect 32030 31220 32036 31232
rect 32088 31220 32094 31272
rect 34054 31220 34060 31272
rect 34112 31260 34118 31272
rect 35345 31263 35403 31269
rect 35345 31260 35357 31263
rect 34112 31232 35357 31260
rect 34112 31220 34118 31232
rect 35345 31229 35357 31232
rect 35391 31229 35403 31263
rect 35345 31223 35403 31229
rect 36725 31195 36783 31201
rect 33428 31164 33916 31192
rect 33428 31124 33456 31164
rect 27540 31096 33456 31124
rect 33505 31127 33563 31133
rect 33505 31093 33517 31127
rect 33551 31124 33563 31127
rect 33778 31124 33784 31136
rect 33551 31096 33784 31124
rect 33551 31093 33563 31096
rect 33505 31087 33563 31093
rect 33778 31084 33784 31096
rect 33836 31084 33842 31136
rect 33888 31124 33916 31164
rect 36725 31161 36737 31195
rect 36771 31192 36783 31195
rect 37734 31192 37740 31204
rect 36771 31164 37740 31192
rect 36771 31161 36783 31164
rect 36725 31155 36783 31161
rect 37734 31152 37740 31164
rect 37792 31152 37798 31204
rect 37550 31124 37556 31136
rect 33888 31096 37556 31124
rect 37550 31084 37556 31096
rect 37608 31084 37614 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 2130 30880 2136 30932
rect 2188 30920 2194 30932
rect 25866 30920 25872 30932
rect 2188 30892 22094 30920
rect 25827 30892 25872 30920
rect 2188 30880 2194 30892
rect 16301 30855 16359 30861
rect 16301 30821 16313 30855
rect 16347 30852 16359 30855
rect 16666 30852 16672 30864
rect 16347 30824 16672 30852
rect 16347 30821 16359 30824
rect 16301 30815 16359 30821
rect 16666 30812 16672 30824
rect 16724 30812 16730 30864
rect 16761 30855 16819 30861
rect 16761 30821 16773 30855
rect 16807 30852 16819 30855
rect 17034 30852 17040 30864
rect 16807 30824 17040 30852
rect 16807 30821 16819 30824
rect 16761 30815 16819 30821
rect 17034 30812 17040 30824
rect 17092 30812 17098 30864
rect 20622 30812 20628 30864
rect 20680 30852 20686 30864
rect 20809 30855 20867 30861
rect 20809 30852 20821 30855
rect 20680 30824 20821 30852
rect 20680 30812 20686 30824
rect 20809 30821 20821 30824
rect 20855 30821 20867 30855
rect 20809 30815 20867 30821
rect 19889 30787 19947 30793
rect 19889 30753 19901 30787
rect 19935 30784 19947 30787
rect 21177 30787 21235 30793
rect 19935 30756 20852 30784
rect 19935 30753 19947 30756
rect 19889 30747 19947 30753
rect 20824 30728 20852 30756
rect 21177 30753 21189 30787
rect 21223 30784 21235 30787
rect 21266 30784 21272 30796
rect 21223 30756 21272 30784
rect 21223 30753 21235 30756
rect 21177 30747 21235 30753
rect 21266 30744 21272 30756
rect 21324 30744 21330 30796
rect 22066 30784 22094 30892
rect 25866 30880 25872 30892
rect 25924 30880 25930 30932
rect 27522 30920 27528 30932
rect 27483 30892 27528 30920
rect 27522 30880 27528 30892
rect 27580 30880 27586 30932
rect 28537 30923 28595 30929
rect 27632 30892 28212 30920
rect 24486 30812 24492 30864
rect 24544 30852 24550 30864
rect 24581 30855 24639 30861
rect 24581 30852 24593 30855
rect 24544 30824 24593 30852
rect 24544 30812 24550 30824
rect 24581 30821 24593 30824
rect 24627 30821 24639 30855
rect 24581 30815 24639 30821
rect 27632 30784 27660 30892
rect 22066 30756 27660 30784
rect 28184 30784 28212 30892
rect 28537 30889 28549 30923
rect 28583 30920 28595 30923
rect 29454 30920 29460 30932
rect 28583 30892 29460 30920
rect 28583 30889 28595 30892
rect 28537 30883 28595 30889
rect 29454 30880 29460 30892
rect 29512 30880 29518 30932
rect 29730 30880 29736 30932
rect 29788 30920 29794 30932
rect 30377 30923 30435 30929
rect 30377 30920 30389 30923
rect 29788 30892 30389 30920
rect 29788 30880 29794 30892
rect 30377 30889 30389 30892
rect 30423 30889 30435 30923
rect 30377 30883 30435 30889
rect 28626 30812 28632 30864
rect 28684 30852 28690 30864
rect 29549 30855 29607 30861
rect 29549 30852 29561 30855
rect 28684 30824 29561 30852
rect 28684 30812 28690 30824
rect 29549 30821 29561 30824
rect 29595 30821 29607 30855
rect 29549 30815 29607 30821
rect 32398 30784 32404 30796
rect 28184 30756 32404 30784
rect 32398 30744 32404 30756
rect 32456 30744 32462 30796
rect 37182 30784 37188 30796
rect 37143 30756 37188 30784
rect 37182 30744 37188 30756
rect 37240 30744 37246 30796
rect 37274 30744 37280 30796
rect 37332 30784 37338 30796
rect 37918 30784 37924 30796
rect 37332 30756 37924 30784
rect 37332 30744 37338 30756
rect 37918 30744 37924 30756
rect 37976 30744 37982 30796
rect 14274 30716 14280 30728
rect 14235 30688 14280 30716
rect 14274 30676 14280 30688
rect 14332 30676 14338 30728
rect 14921 30719 14979 30725
rect 14921 30685 14933 30719
rect 14967 30716 14979 30719
rect 18046 30716 18052 30728
rect 14967 30688 18052 30716
rect 14967 30685 14979 30688
rect 14921 30679 14979 30685
rect 18046 30676 18052 30688
rect 18104 30716 18110 30728
rect 18141 30719 18199 30725
rect 18141 30716 18153 30719
rect 18104 30688 18153 30716
rect 18104 30676 18110 30688
rect 18141 30685 18153 30688
rect 18187 30716 18199 30719
rect 18414 30716 18420 30728
rect 18187 30688 18420 30716
rect 18187 30685 18199 30688
rect 18141 30679 18199 30685
rect 18414 30676 18420 30688
rect 18472 30676 18478 30728
rect 20070 30716 20076 30728
rect 20031 30688 20076 30716
rect 20070 30676 20076 30688
rect 20128 30676 20134 30728
rect 20806 30676 20812 30728
rect 20864 30716 20870 30728
rect 21637 30719 21695 30725
rect 21637 30716 21649 30719
rect 20864 30688 21649 30716
rect 20864 30676 20870 30688
rect 21637 30685 21649 30688
rect 21683 30685 21695 30719
rect 21818 30716 21824 30728
rect 21779 30688 21824 30716
rect 21637 30679 21695 30685
rect 21818 30676 21824 30688
rect 21876 30676 21882 30728
rect 22830 30676 22836 30728
rect 22888 30716 22894 30728
rect 23017 30719 23075 30725
rect 23017 30716 23029 30719
rect 22888 30688 23029 30716
rect 22888 30676 22894 30688
rect 23017 30685 23029 30688
rect 23063 30685 23075 30719
rect 24762 30716 24768 30728
rect 24723 30688 24768 30716
rect 23017 30679 23075 30685
rect 24762 30676 24768 30688
rect 24820 30676 24826 30728
rect 25317 30719 25375 30725
rect 25317 30685 25329 30719
rect 25363 30685 25375 30719
rect 25498 30716 25504 30728
rect 25459 30688 25504 30716
rect 25317 30679 25375 30685
rect 15166 30651 15224 30657
rect 15166 30648 15178 30651
rect 14476 30620 15178 30648
rect 14476 30589 14504 30620
rect 15166 30617 15178 30620
rect 15212 30617 15224 30651
rect 15166 30611 15224 30617
rect 17678 30608 17684 30660
rect 17736 30648 17742 30660
rect 17874 30651 17932 30657
rect 17874 30648 17886 30651
rect 17736 30620 17886 30648
rect 17736 30608 17742 30620
rect 17874 30617 17886 30620
rect 17920 30617 17932 30651
rect 17874 30611 17932 30617
rect 20257 30651 20315 30657
rect 20257 30617 20269 30651
rect 20303 30648 20315 30651
rect 20898 30648 20904 30660
rect 20303 30620 20904 30648
rect 20303 30617 20315 30620
rect 20257 30611 20315 30617
rect 20898 30608 20904 30620
rect 20956 30608 20962 30660
rect 24486 30608 24492 30660
rect 24544 30648 24550 30660
rect 25332 30648 25360 30679
rect 25498 30676 25504 30688
rect 25556 30676 25562 30728
rect 25685 30719 25743 30725
rect 25685 30685 25697 30719
rect 25731 30716 25743 30719
rect 26970 30716 26976 30728
rect 25731 30688 26976 30716
rect 25731 30685 25743 30688
rect 25685 30679 25743 30685
rect 26970 30676 26976 30688
rect 27028 30716 27034 30728
rect 27249 30719 27307 30725
rect 27249 30716 27261 30719
rect 27028 30688 27261 30716
rect 27028 30676 27034 30688
rect 27249 30685 27261 30688
rect 27295 30685 27307 30719
rect 27249 30679 27307 30685
rect 27341 30719 27399 30725
rect 27341 30685 27353 30719
rect 27387 30685 27399 30719
rect 27341 30679 27399 30685
rect 24544 30620 25360 30648
rect 25593 30651 25651 30657
rect 24544 30608 24550 30620
rect 25593 30617 25605 30651
rect 25639 30648 25651 30651
rect 26418 30648 26424 30660
rect 25639 30620 26424 30648
rect 25639 30617 25651 30620
rect 25593 30611 25651 30617
rect 26418 30608 26424 30620
rect 26476 30648 26482 30660
rect 27356 30648 27384 30679
rect 27430 30676 27436 30728
rect 27488 30716 27494 30728
rect 27617 30719 27675 30725
rect 27617 30716 27629 30719
rect 27488 30688 27629 30716
rect 27488 30676 27494 30688
rect 27617 30685 27629 30688
rect 27663 30685 27675 30719
rect 28074 30716 28080 30728
rect 28035 30688 28080 30716
rect 27617 30679 27675 30685
rect 26476 30620 27384 30648
rect 27632 30648 27660 30679
rect 28074 30676 28080 30688
rect 28132 30676 28138 30728
rect 28350 30716 28356 30728
rect 28311 30688 28356 30716
rect 28350 30676 28356 30688
rect 28408 30676 28414 30728
rect 30469 30719 30527 30725
rect 30469 30685 30481 30719
rect 30515 30716 30527 30719
rect 30926 30716 30932 30728
rect 30515 30688 30932 30716
rect 30515 30685 30527 30688
rect 30469 30679 30527 30685
rect 30926 30676 30932 30688
rect 30984 30676 30990 30728
rect 31846 30716 31852 30728
rect 31807 30688 31852 30716
rect 31846 30676 31852 30688
rect 31904 30676 31910 30728
rect 38105 30719 38163 30725
rect 38105 30685 38117 30719
rect 38151 30716 38163 30719
rect 38194 30716 38200 30728
rect 38151 30688 38200 30716
rect 38151 30685 38163 30688
rect 38105 30679 38163 30685
rect 38194 30676 38200 30688
rect 38252 30676 38258 30728
rect 29733 30651 29791 30657
rect 29733 30648 29745 30651
rect 27632 30620 29745 30648
rect 26476 30608 26482 30620
rect 29733 30617 29745 30620
rect 29779 30617 29791 30651
rect 37918 30648 37924 30660
rect 37879 30620 37924 30648
rect 29733 30611 29791 30617
rect 37918 30608 37924 30620
rect 37976 30608 37982 30660
rect 14461 30583 14519 30589
rect 14461 30549 14473 30583
rect 14507 30549 14519 30583
rect 14461 30543 14519 30549
rect 20717 30583 20775 30589
rect 20717 30549 20729 30583
rect 20763 30580 20775 30583
rect 21082 30580 21088 30592
rect 20763 30552 21088 30580
rect 20763 30549 20775 30552
rect 20717 30543 20775 30549
rect 21082 30540 21088 30552
rect 21140 30540 21146 30592
rect 21729 30583 21787 30589
rect 21729 30549 21741 30583
rect 21775 30580 21787 30583
rect 21910 30580 21916 30592
rect 21775 30552 21916 30580
rect 21775 30549 21787 30552
rect 21729 30543 21787 30549
rect 21910 30540 21916 30552
rect 21968 30540 21974 30592
rect 23201 30583 23259 30589
rect 23201 30549 23213 30583
rect 23247 30580 23259 30583
rect 23290 30580 23296 30592
rect 23247 30552 23296 30580
rect 23247 30549 23259 30552
rect 23201 30543 23259 30549
rect 23290 30540 23296 30552
rect 23348 30580 23354 30592
rect 26602 30580 26608 30592
rect 23348 30552 26608 30580
rect 23348 30540 23354 30552
rect 26602 30540 26608 30552
rect 26660 30540 26666 30592
rect 27065 30583 27123 30589
rect 27065 30549 27077 30583
rect 27111 30580 27123 30583
rect 28169 30583 28227 30589
rect 28169 30580 28181 30583
rect 27111 30552 28181 30580
rect 27111 30549 27123 30552
rect 27065 30543 27123 30549
rect 28169 30549 28181 30552
rect 28215 30549 28227 30583
rect 28169 30543 28227 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 21082 30336 21088 30388
rect 21140 30376 21146 30388
rect 22002 30376 22008 30388
rect 21140 30348 22008 30376
rect 21140 30336 21146 30348
rect 22002 30336 22008 30348
rect 22060 30336 22066 30388
rect 27522 30376 27528 30388
rect 27483 30348 27528 30376
rect 27522 30336 27528 30348
rect 27580 30336 27586 30388
rect 28736 30348 29040 30376
rect 24949 30311 25007 30317
rect 15396 30280 24532 30308
rect 14918 30240 14924 30252
rect 14879 30212 14924 30240
rect 14918 30200 14924 30212
rect 14976 30200 14982 30252
rect 15396 30184 15424 30280
rect 18598 30240 18604 30252
rect 18559 30212 18604 30240
rect 18598 30200 18604 30212
rect 18656 30200 18662 30252
rect 20533 30243 20591 30249
rect 20533 30209 20545 30243
rect 20579 30209 20591 30243
rect 20533 30203 20591 30209
rect 20717 30243 20775 30249
rect 20717 30209 20729 30243
rect 20763 30209 20775 30243
rect 20898 30240 20904 30252
rect 20859 30212 20904 30240
rect 20717 30203 20775 30209
rect 15378 30172 15384 30184
rect 15339 30144 15384 30172
rect 15378 30132 15384 30144
rect 15436 30132 15442 30184
rect 18417 30039 18475 30045
rect 18417 30005 18429 30039
rect 18463 30036 18475 30039
rect 18598 30036 18604 30048
rect 18463 30008 18604 30036
rect 18463 30005 18475 30008
rect 18417 29999 18475 30005
rect 18598 29996 18604 30008
rect 18656 29996 18662 30048
rect 20548 30036 20576 30203
rect 20732 30104 20760 30203
rect 20898 30200 20904 30212
rect 20956 30200 20962 30252
rect 21082 30240 21088 30252
rect 21043 30212 21088 30240
rect 21082 30200 21088 30212
rect 21140 30200 21146 30252
rect 21542 30200 21548 30252
rect 21600 30240 21606 30252
rect 21910 30240 21916 30252
rect 21600 30212 21916 30240
rect 21600 30200 21606 30212
rect 21910 30200 21916 30212
rect 21968 30240 21974 30252
rect 22005 30243 22063 30249
rect 22005 30240 22017 30243
rect 21968 30212 22017 30240
rect 21968 30200 21974 30212
rect 22005 30209 22017 30212
rect 22051 30209 22063 30243
rect 22005 30203 22063 30209
rect 22094 30200 22100 30252
rect 22152 30240 22158 30252
rect 22281 30243 22339 30249
rect 22152 30212 22197 30240
rect 22152 30200 22158 30212
rect 22281 30209 22293 30243
rect 22327 30209 22339 30243
rect 22281 30203 22339 30209
rect 20809 30175 20867 30181
rect 20809 30141 20821 30175
rect 20855 30172 20867 30175
rect 20990 30172 20996 30184
rect 20855 30144 20996 30172
rect 20855 30141 20867 30144
rect 20809 30135 20867 30141
rect 20990 30132 20996 30144
rect 21048 30132 21054 30184
rect 21174 30132 21180 30184
rect 21232 30172 21238 30184
rect 22186 30172 22192 30184
rect 21232 30144 22192 30172
rect 21232 30132 21238 30144
rect 22186 30132 22192 30144
rect 22244 30172 22250 30184
rect 22296 30172 22324 30203
rect 22370 30200 22376 30252
rect 22428 30240 22434 30252
rect 22428 30212 22473 30240
rect 22428 30200 22434 30212
rect 22244 30144 22324 30172
rect 24504 30172 24532 30280
rect 24949 30277 24961 30311
rect 24995 30308 25007 30311
rect 26326 30308 26332 30320
rect 24995 30280 26332 30308
rect 24995 30277 25007 30280
rect 24949 30271 25007 30277
rect 26326 30268 26332 30280
rect 26384 30268 26390 30320
rect 28736 30308 28764 30348
rect 28902 30308 28908 30320
rect 28368 30280 28764 30308
rect 28863 30280 28908 30308
rect 24578 30200 24584 30252
rect 24636 30240 24642 30252
rect 24857 30243 24915 30249
rect 24857 30240 24869 30243
rect 24636 30212 24869 30240
rect 24636 30200 24642 30212
rect 24857 30209 24869 30212
rect 24903 30209 24915 30243
rect 25038 30240 25044 30252
rect 24999 30212 25044 30240
rect 24857 30203 24915 30209
rect 25038 30200 25044 30212
rect 25096 30200 25102 30252
rect 27617 30243 27675 30249
rect 27617 30209 27629 30243
rect 27663 30240 27675 30243
rect 28258 30240 28264 30252
rect 27663 30212 28264 30240
rect 27663 30209 27675 30212
rect 27617 30203 27675 30209
rect 28258 30200 28264 30212
rect 28316 30200 28322 30252
rect 28368 30249 28396 30280
rect 28902 30268 28908 30280
rect 28960 30268 28966 30320
rect 29012 30308 29040 30348
rect 30392 30348 30696 30376
rect 30392 30308 30420 30348
rect 29012 30280 30420 30308
rect 30460 30311 30518 30317
rect 30460 30277 30472 30311
rect 30506 30308 30518 30311
rect 30558 30308 30564 30320
rect 30506 30280 30564 30308
rect 30506 30277 30518 30280
rect 30460 30271 30518 30277
rect 30558 30268 30564 30280
rect 30616 30268 30622 30320
rect 30668 30308 30696 30348
rect 31294 30336 31300 30388
rect 31352 30376 31358 30388
rect 31573 30379 31631 30385
rect 31573 30376 31585 30379
rect 31352 30348 31585 30376
rect 31352 30336 31358 30348
rect 31573 30345 31585 30348
rect 31619 30345 31631 30379
rect 31573 30339 31631 30345
rect 37461 30379 37519 30385
rect 37461 30345 37473 30379
rect 37507 30376 37519 30379
rect 37918 30376 37924 30388
rect 37507 30348 37924 30376
rect 37507 30345 37519 30348
rect 37461 30339 37519 30345
rect 37918 30336 37924 30348
rect 37976 30336 37982 30388
rect 31478 30308 31484 30320
rect 30668 30280 31484 30308
rect 31478 30268 31484 30280
rect 31536 30268 31542 30320
rect 33137 30311 33195 30317
rect 33137 30277 33149 30311
rect 33183 30308 33195 30311
rect 33318 30308 33324 30320
rect 33183 30280 33324 30308
rect 33183 30277 33195 30280
rect 33137 30271 33195 30277
rect 33318 30268 33324 30280
rect 33376 30268 33382 30320
rect 34324 30311 34382 30317
rect 34324 30277 34336 30311
rect 34370 30308 34382 30311
rect 34422 30308 34428 30320
rect 34370 30280 34428 30308
rect 34370 30277 34382 30280
rect 34324 30271 34382 30277
rect 34422 30268 34428 30280
rect 34480 30268 34486 30320
rect 28353 30243 28411 30249
rect 28353 30209 28365 30243
rect 28399 30209 28411 30243
rect 28810 30240 28816 30252
rect 28771 30212 28816 30240
rect 28353 30203 28411 30209
rect 28810 30200 28816 30212
rect 28868 30200 28874 30252
rect 28994 30200 29000 30252
rect 29052 30240 29058 30252
rect 29457 30243 29515 30249
rect 29457 30240 29469 30243
rect 29052 30212 29469 30240
rect 29052 30200 29058 30212
rect 29457 30209 29469 30212
rect 29503 30209 29515 30243
rect 29638 30240 29644 30252
rect 29599 30212 29644 30240
rect 29457 30203 29515 30209
rect 29638 30200 29644 30212
rect 29696 30200 29702 30252
rect 34054 30240 34060 30252
rect 29748 30212 31754 30240
rect 34015 30212 34060 30240
rect 29748 30172 29776 30212
rect 24504 30144 29776 30172
rect 30193 30175 30251 30181
rect 22244 30132 22250 30144
rect 30193 30141 30205 30175
rect 30239 30141 30251 30175
rect 31726 30172 31754 30212
rect 34054 30200 34060 30212
rect 34112 30200 34118 30252
rect 37274 30240 37280 30252
rect 34164 30212 37280 30240
rect 34164 30172 34192 30212
rect 37274 30200 37280 30212
rect 37332 30200 37338 30252
rect 37369 30243 37427 30249
rect 37369 30209 37381 30243
rect 37415 30240 37427 30243
rect 37458 30240 37464 30252
rect 37415 30212 37464 30240
rect 37415 30209 37427 30212
rect 37369 30203 37427 30209
rect 37458 30200 37464 30212
rect 37516 30200 37522 30252
rect 31726 30144 34192 30172
rect 30193 30135 30251 30141
rect 20898 30104 20904 30116
rect 20732 30076 20904 30104
rect 20898 30064 20904 30076
rect 20956 30064 20962 30116
rect 21358 30104 21364 30116
rect 21100 30076 21364 30104
rect 21100 30036 21128 30076
rect 21358 30064 21364 30076
rect 21416 30064 21422 30116
rect 27890 30064 27896 30116
rect 27948 30104 27954 30116
rect 28169 30107 28227 30113
rect 28169 30104 28181 30107
rect 27948 30076 28181 30104
rect 27948 30064 27954 30076
rect 28169 30073 28181 30076
rect 28215 30073 28227 30107
rect 28169 30067 28227 30073
rect 21266 30036 21272 30048
rect 20548 30008 21128 30036
rect 21227 30008 21272 30036
rect 21266 29996 21272 30008
rect 21324 29996 21330 30048
rect 21818 30036 21824 30048
rect 21779 30008 21824 30036
rect 21818 29996 21824 30008
rect 21876 29996 21882 30048
rect 29454 30036 29460 30048
rect 29415 30008 29460 30036
rect 29454 29996 29460 30008
rect 29512 29996 29518 30048
rect 30208 30036 30236 30135
rect 31570 30064 31576 30116
rect 31628 30104 31634 30116
rect 31754 30104 31760 30116
rect 31628 30076 31760 30104
rect 31628 30064 31634 30076
rect 31754 30064 31760 30076
rect 31812 30064 31818 30116
rect 33226 30064 33232 30116
rect 33284 30104 33290 30116
rect 33413 30107 33471 30113
rect 33413 30104 33425 30107
rect 33284 30076 33425 30104
rect 33284 30064 33290 30076
rect 33413 30073 33425 30076
rect 33459 30073 33471 30107
rect 33413 30067 33471 30073
rect 30374 30036 30380 30048
rect 30208 30008 30380 30036
rect 30374 29996 30380 30008
rect 30432 30036 30438 30048
rect 31662 30036 31668 30048
rect 30432 30008 31668 30036
rect 30432 29996 30438 30008
rect 31662 29996 31668 30008
rect 31720 29996 31726 30048
rect 33597 30039 33655 30045
rect 33597 30005 33609 30039
rect 33643 30036 33655 30039
rect 33686 30036 33692 30048
rect 33643 30008 33692 30036
rect 33643 30005 33655 30008
rect 33597 29999 33655 30005
rect 33686 29996 33692 30008
rect 33744 29996 33750 30048
rect 35434 30036 35440 30048
rect 35395 30008 35440 30036
rect 35434 29996 35440 30008
rect 35492 29996 35498 30048
rect 36262 29996 36268 30048
rect 36320 30036 36326 30048
rect 36541 30039 36599 30045
rect 36541 30036 36553 30039
rect 36320 30008 36553 30036
rect 36320 29996 36326 30008
rect 36541 30005 36553 30008
rect 36587 30005 36599 30039
rect 36541 29999 36599 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 20990 29792 20996 29844
rect 21048 29832 21054 29844
rect 21085 29835 21143 29841
rect 21085 29832 21097 29835
rect 21048 29804 21097 29832
rect 21048 29792 21054 29804
rect 21085 29801 21097 29804
rect 21131 29801 21143 29835
rect 25409 29835 25467 29841
rect 21085 29795 21143 29801
rect 21192 29804 25360 29832
rect 15654 29696 15660 29708
rect 15615 29668 15660 29696
rect 15654 29656 15660 29668
rect 15712 29656 15718 29708
rect 18598 29656 18604 29708
rect 18656 29696 18662 29708
rect 21192 29696 21220 29804
rect 21358 29724 21364 29776
rect 21416 29764 21422 29776
rect 22370 29764 22376 29776
rect 21416 29736 22376 29764
rect 21416 29724 21422 29736
rect 22370 29724 22376 29736
rect 22428 29764 22434 29776
rect 22830 29764 22836 29776
rect 22428 29736 22836 29764
rect 22428 29724 22434 29736
rect 22830 29724 22836 29736
rect 22888 29724 22894 29776
rect 21634 29696 21640 29708
rect 18656 29668 21220 29696
rect 21595 29668 21640 29696
rect 18656 29656 18662 29668
rect 21634 29656 21640 29668
rect 21692 29656 21698 29708
rect 22186 29696 22192 29708
rect 21836 29668 22192 29696
rect 1670 29588 1676 29640
rect 1728 29628 1734 29640
rect 1765 29631 1823 29637
rect 1765 29628 1777 29631
rect 1728 29600 1777 29628
rect 1728 29588 1734 29600
rect 1765 29597 1777 29600
rect 1811 29597 1823 29631
rect 14182 29628 14188 29640
rect 14143 29600 14188 29628
rect 1765 29591 1823 29597
rect 14182 29588 14188 29600
rect 14240 29588 14246 29640
rect 14918 29588 14924 29640
rect 14976 29628 14982 29640
rect 15289 29631 15347 29637
rect 15289 29628 15301 29631
rect 14976 29600 15301 29628
rect 14976 29588 14982 29600
rect 15289 29597 15301 29600
rect 15335 29597 15347 29631
rect 20806 29628 20812 29640
rect 20767 29600 20812 29628
rect 15289 29591 15347 29597
rect 20806 29588 20812 29600
rect 20864 29588 20870 29640
rect 20898 29588 20904 29640
rect 20956 29628 20962 29640
rect 20956 29600 21049 29628
rect 20956 29588 20962 29600
rect 21082 29588 21088 29640
rect 21140 29628 21146 29640
rect 21836 29637 21864 29668
rect 22186 29656 22192 29668
rect 22244 29656 22250 29708
rect 25332 29696 25360 29804
rect 25409 29801 25421 29835
rect 25455 29832 25467 29835
rect 25498 29832 25504 29844
rect 25455 29804 25504 29832
rect 25455 29801 25467 29804
rect 25409 29795 25467 29801
rect 25498 29792 25504 29804
rect 25556 29792 25562 29844
rect 26050 29832 26056 29844
rect 26011 29804 26056 29832
rect 26050 29792 26056 29804
rect 26108 29792 26114 29844
rect 26970 29832 26976 29844
rect 26931 29804 26976 29832
rect 26970 29792 26976 29804
rect 27028 29792 27034 29844
rect 28813 29835 28871 29841
rect 28813 29801 28825 29835
rect 28859 29832 28871 29835
rect 28994 29832 29000 29844
rect 28859 29804 29000 29832
rect 28859 29801 28871 29804
rect 28813 29795 28871 29801
rect 28994 29792 29000 29804
rect 29052 29792 29058 29844
rect 30926 29832 30932 29844
rect 29472 29804 30932 29832
rect 27154 29696 27160 29708
rect 25332 29668 27160 29696
rect 27154 29656 27160 29668
rect 27212 29696 27218 29708
rect 28721 29699 28779 29705
rect 28721 29696 28733 29699
rect 27212 29668 28733 29696
rect 27212 29656 27218 29668
rect 28721 29665 28733 29668
rect 28767 29665 28779 29699
rect 28721 29659 28779 29665
rect 21177 29631 21235 29637
rect 21177 29628 21189 29631
rect 21140 29600 21189 29628
rect 21140 29588 21146 29600
rect 21177 29597 21189 29600
rect 21223 29597 21235 29631
rect 21177 29591 21235 29597
rect 21821 29631 21879 29637
rect 21821 29597 21833 29631
rect 21867 29597 21879 29631
rect 22002 29628 22008 29640
rect 21963 29600 22008 29628
rect 21821 29591 21879 29597
rect 22002 29588 22008 29600
rect 22060 29588 22066 29640
rect 22097 29631 22155 29637
rect 22097 29597 22109 29631
rect 22143 29597 22155 29631
rect 23106 29628 23112 29640
rect 23067 29600 23112 29628
rect 22097 29591 22155 29597
rect 15654 29520 15660 29572
rect 15712 29560 15718 29572
rect 20916 29560 20944 29588
rect 21542 29560 21548 29572
rect 15712 29532 20852 29560
rect 20916 29532 21548 29560
rect 15712 29520 15718 29532
rect 14366 29492 14372 29504
rect 14327 29464 14372 29492
rect 14366 29452 14372 29464
rect 14424 29452 14430 29504
rect 20622 29492 20628 29504
rect 20583 29464 20628 29492
rect 20622 29452 20628 29464
rect 20680 29452 20686 29504
rect 20824 29492 20852 29532
rect 21542 29520 21548 29532
rect 21600 29560 21606 29572
rect 22112 29560 22140 29591
rect 23106 29588 23112 29600
rect 23164 29588 23170 29640
rect 25498 29628 25504 29640
rect 25459 29600 25504 29628
rect 25498 29588 25504 29600
rect 25556 29588 25562 29640
rect 25958 29628 25964 29640
rect 25919 29600 25964 29628
rect 25958 29588 25964 29600
rect 26016 29588 26022 29640
rect 26878 29628 26884 29640
rect 26839 29600 26884 29628
rect 26878 29588 26884 29600
rect 26936 29588 26942 29640
rect 28902 29628 28908 29640
rect 28863 29600 28908 29628
rect 28902 29588 28908 29600
rect 28960 29588 28966 29640
rect 28997 29631 29055 29637
rect 28997 29597 29009 29631
rect 29043 29628 29055 29631
rect 29270 29628 29276 29640
rect 29043 29600 29276 29628
rect 29043 29597 29055 29600
rect 28997 29591 29055 29597
rect 29270 29588 29276 29600
rect 29328 29628 29334 29640
rect 29472 29628 29500 29804
rect 30926 29792 30932 29804
rect 30984 29792 30990 29844
rect 30650 29724 30656 29776
rect 30708 29764 30714 29776
rect 31389 29767 31447 29773
rect 31389 29764 31401 29767
rect 30708 29736 31401 29764
rect 30708 29724 30714 29736
rect 31389 29733 31401 29736
rect 31435 29733 31447 29767
rect 31389 29727 31447 29733
rect 32953 29767 33011 29773
rect 32953 29733 32965 29767
rect 32999 29764 33011 29767
rect 33318 29764 33324 29776
rect 32999 29736 33324 29764
rect 32999 29733 33011 29736
rect 32953 29727 33011 29733
rect 33318 29724 33324 29736
rect 33376 29764 33382 29776
rect 34149 29767 34207 29773
rect 33376 29736 33548 29764
rect 33376 29724 33382 29736
rect 33520 29705 33548 29736
rect 34149 29733 34161 29767
rect 34195 29764 34207 29767
rect 34790 29764 34796 29776
rect 34195 29736 34796 29764
rect 34195 29733 34207 29736
rect 34149 29727 34207 29733
rect 34790 29724 34796 29736
rect 34848 29724 34854 29776
rect 33505 29699 33563 29705
rect 33505 29665 33517 29699
rect 33551 29665 33563 29699
rect 33778 29696 33784 29708
rect 33739 29668 33784 29696
rect 33505 29659 33563 29665
rect 33778 29656 33784 29668
rect 33836 29656 33842 29708
rect 35434 29696 35440 29708
rect 34900 29668 35440 29696
rect 29328 29600 29500 29628
rect 29549 29631 29607 29637
rect 29328 29588 29334 29600
rect 29549 29597 29561 29631
rect 29595 29628 29607 29631
rect 30374 29628 30380 29640
rect 29595 29600 30380 29628
rect 29595 29597 29607 29600
rect 29549 29591 29607 29597
rect 30374 29588 30380 29600
rect 30432 29588 30438 29640
rect 31662 29628 31668 29640
rect 31623 29600 31668 29628
rect 31662 29588 31668 29600
rect 31720 29588 31726 29640
rect 33873 29631 33931 29637
rect 33873 29597 33885 29631
rect 33919 29628 33931 29631
rect 34606 29628 34612 29640
rect 33919 29600 34612 29628
rect 33919 29597 33931 29600
rect 33873 29591 33931 29597
rect 34606 29588 34612 29600
rect 34664 29628 34670 29640
rect 34900 29637 34928 29668
rect 35434 29656 35440 29668
rect 35492 29656 35498 29708
rect 36262 29696 36268 29708
rect 36223 29668 36268 29696
rect 36262 29656 36268 29668
rect 36320 29656 36326 29708
rect 38102 29696 38108 29708
rect 38063 29668 38108 29696
rect 38102 29656 38108 29668
rect 38160 29656 38166 29708
rect 34885 29631 34943 29637
rect 34885 29628 34897 29631
rect 34664 29600 34897 29628
rect 34664 29588 34670 29600
rect 34885 29597 34897 29600
rect 34931 29597 34943 29631
rect 34885 29591 34943 29597
rect 34977 29631 35035 29637
rect 34977 29597 34989 29631
rect 35023 29597 35035 29631
rect 34977 29591 35035 29597
rect 29362 29560 29368 29572
rect 21600 29532 22140 29560
rect 23124 29532 29368 29560
rect 21600 29520 21606 29532
rect 23124 29492 23152 29532
rect 29362 29520 29368 29532
rect 29420 29520 29426 29572
rect 29454 29520 29460 29572
rect 29512 29560 29518 29572
rect 29794 29563 29852 29569
rect 29794 29560 29806 29563
rect 29512 29532 29806 29560
rect 29512 29520 29518 29532
rect 29794 29529 29806 29532
rect 29840 29529 29852 29563
rect 29794 29523 29852 29529
rect 30834 29520 30840 29572
rect 30892 29560 30898 29572
rect 31389 29563 31447 29569
rect 31389 29560 31401 29563
rect 30892 29532 31401 29560
rect 30892 29520 30898 29532
rect 31389 29529 31401 29532
rect 31435 29529 31447 29563
rect 31389 29523 31447 29529
rect 32585 29563 32643 29569
rect 32585 29529 32597 29563
rect 32631 29560 32643 29563
rect 33226 29560 33232 29572
rect 32631 29532 33232 29560
rect 32631 29529 32643 29532
rect 32585 29523 32643 29529
rect 33226 29520 33232 29532
rect 33284 29560 33290 29572
rect 33990 29563 34048 29569
rect 33990 29560 34002 29563
rect 33284 29532 34002 29560
rect 33284 29520 33290 29532
rect 33990 29529 34002 29532
rect 34036 29529 34048 29563
rect 33990 29523 34048 29529
rect 34422 29520 34428 29572
rect 34480 29560 34486 29572
rect 34992 29560 35020 29591
rect 34480 29532 35020 29560
rect 36449 29563 36507 29569
rect 34480 29520 34486 29532
rect 36449 29529 36461 29563
rect 36495 29560 36507 29563
rect 37366 29560 37372 29572
rect 36495 29532 37372 29560
rect 36495 29529 36507 29532
rect 36449 29523 36507 29529
rect 37366 29520 37372 29532
rect 37424 29520 37430 29572
rect 23290 29492 23296 29504
rect 20824 29464 23152 29492
rect 23251 29464 23296 29492
rect 23290 29452 23296 29464
rect 23348 29452 23354 29504
rect 24854 29452 24860 29504
rect 24912 29492 24918 29504
rect 31202 29492 31208 29504
rect 24912 29464 31208 29492
rect 24912 29452 24918 29464
rect 31202 29452 31208 29464
rect 31260 29452 31266 29504
rect 31294 29452 31300 29504
rect 31352 29492 31358 29504
rect 31573 29495 31631 29501
rect 31573 29492 31585 29495
rect 31352 29464 31585 29492
rect 31352 29452 31358 29464
rect 31573 29461 31585 29464
rect 31619 29461 31631 29495
rect 31573 29455 31631 29461
rect 33045 29495 33103 29501
rect 33045 29461 33057 29495
rect 33091 29492 33103 29495
rect 33410 29492 33416 29504
rect 33091 29464 33416 29492
rect 33091 29461 33103 29464
rect 33045 29455 33103 29461
rect 33410 29452 33416 29464
rect 33468 29452 33474 29504
rect 34514 29452 34520 29504
rect 34572 29492 34578 29504
rect 34701 29495 34759 29501
rect 34701 29492 34713 29495
rect 34572 29464 34713 29492
rect 34572 29452 34578 29464
rect 34701 29461 34713 29464
rect 34747 29461 34759 29495
rect 34701 29455 34759 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 24854 29288 24860 29300
rect 14384 29260 24860 29288
rect 14384 29220 14412 29260
rect 24854 29248 24860 29260
rect 24912 29248 24918 29300
rect 24949 29291 25007 29297
rect 24949 29257 24961 29291
rect 24995 29288 25007 29291
rect 25406 29288 25412 29300
rect 24995 29260 25412 29288
rect 24995 29257 25007 29260
rect 24949 29251 25007 29257
rect 25406 29248 25412 29260
rect 25464 29288 25470 29300
rect 25958 29288 25964 29300
rect 25464 29260 25964 29288
rect 25464 29248 25470 29260
rect 25958 29248 25964 29260
rect 26016 29248 26022 29300
rect 26878 29248 26884 29300
rect 26936 29288 26942 29300
rect 26973 29291 27031 29297
rect 26973 29288 26985 29291
rect 26936 29260 26985 29288
rect 26936 29248 26942 29260
rect 26973 29257 26985 29260
rect 27019 29257 27031 29291
rect 29638 29288 29644 29300
rect 29599 29260 29644 29288
rect 26973 29251 27031 29257
rect 29638 29248 29644 29260
rect 29696 29248 29702 29300
rect 30469 29291 30527 29297
rect 30469 29257 30481 29291
rect 30515 29288 30527 29291
rect 30558 29288 30564 29300
rect 30515 29260 30564 29288
rect 30515 29257 30527 29260
rect 30469 29251 30527 29257
rect 30558 29248 30564 29260
rect 30616 29248 30622 29300
rect 31662 29288 31668 29300
rect 30852 29260 31668 29288
rect 25133 29223 25191 29229
rect 14200 29192 14412 29220
rect 15672 29192 24808 29220
rect 1670 29152 1676 29164
rect 1631 29124 1676 29152
rect 1670 29112 1676 29124
rect 1728 29112 1734 29164
rect 14090 29152 14096 29164
rect 14003 29124 14096 29152
rect 14090 29112 14096 29124
rect 14148 29152 14154 29164
rect 14200 29152 14228 29192
rect 14366 29152 14372 29164
rect 14148 29124 14228 29152
rect 14279 29124 14372 29152
rect 14148 29112 14154 29124
rect 14366 29112 14372 29124
rect 14424 29152 14430 29164
rect 14918 29152 14924 29164
rect 14424 29124 14924 29152
rect 14424 29112 14430 29124
rect 14918 29112 14924 29124
rect 14976 29112 14982 29164
rect 15672 29096 15700 29192
rect 17957 29155 18015 29161
rect 17957 29121 17969 29155
rect 18003 29152 18015 29155
rect 18046 29152 18052 29164
rect 18003 29124 18052 29152
rect 18003 29121 18015 29124
rect 17957 29115 18015 29121
rect 18046 29112 18052 29124
rect 18104 29112 18110 29164
rect 18230 29161 18236 29164
rect 18224 29115 18236 29161
rect 18288 29152 18294 29164
rect 22462 29152 22468 29164
rect 18288 29124 18324 29152
rect 22066 29124 22468 29152
rect 18230 29112 18236 29115
rect 18288 29112 18294 29124
rect 1854 29084 1860 29096
rect 1815 29056 1860 29084
rect 1854 29044 1860 29056
rect 1912 29044 1918 29096
rect 2774 29084 2780 29096
rect 2735 29056 2780 29084
rect 2774 29044 2780 29056
rect 2832 29044 2838 29096
rect 15654 29084 15660 29096
rect 15615 29056 15660 29084
rect 15654 29044 15660 29056
rect 15712 29044 15718 29096
rect 19337 29019 19395 29025
rect 19337 29006 19349 29019
rect 19383 29006 19395 29019
rect 19334 28994 19340 29006
rect 18138 28908 18144 28960
rect 18196 28948 18202 28960
rect 19306 28954 19340 28994
rect 19392 28954 19398 29006
rect 19306 28948 19334 28954
rect 18196 28920 19334 28948
rect 18196 28908 18202 28920
rect 19426 28908 19432 28960
rect 19484 28948 19490 28960
rect 22066 28948 22094 29124
rect 22462 29112 22468 29124
rect 22520 29112 22526 29164
rect 22738 29161 22744 29164
rect 22732 29115 22744 29161
rect 22796 29152 22802 29164
rect 22796 29124 22832 29152
rect 22738 29112 22744 29115
rect 22796 29112 22802 29124
rect 24780 29084 24808 29192
rect 25133 29189 25145 29223
rect 25179 29220 25191 29223
rect 25498 29220 25504 29232
rect 25179 29192 25504 29220
rect 25179 29189 25191 29192
rect 25133 29183 25191 29189
rect 25498 29180 25504 29192
rect 25556 29180 25562 29232
rect 28718 29220 28724 29232
rect 25608 29192 28724 29220
rect 24857 29155 24915 29161
rect 24857 29121 24869 29155
rect 24903 29152 24915 29155
rect 25314 29152 25320 29164
rect 24903 29124 25320 29152
rect 24903 29121 24915 29124
rect 24857 29115 24915 29121
rect 25314 29112 25320 29124
rect 25372 29112 25378 29164
rect 25608 29084 25636 29192
rect 28718 29180 28724 29192
rect 28776 29180 28782 29232
rect 28902 29180 28908 29232
rect 28960 29220 28966 29232
rect 29656 29220 29684 29248
rect 30852 29220 30880 29260
rect 31662 29248 31668 29260
rect 31720 29248 31726 29300
rect 37366 29288 37372 29300
rect 37327 29260 37372 29288
rect 37366 29248 37372 29260
rect 37424 29248 37430 29300
rect 28960 29192 29500 29220
rect 29656 29192 30880 29220
rect 28960 29180 28966 29192
rect 27614 29112 27620 29164
rect 27672 29152 27678 29164
rect 29472 29161 29500 29192
rect 28086 29155 28144 29161
rect 28086 29152 28098 29155
rect 27672 29124 28098 29152
rect 27672 29112 27678 29124
rect 28086 29121 28098 29124
rect 28132 29121 28144 29155
rect 28086 29115 28144 29121
rect 28353 29155 28411 29161
rect 28353 29121 28365 29155
rect 28399 29121 28411 29155
rect 28353 29115 28411 29121
rect 29457 29155 29515 29161
rect 29457 29121 29469 29155
rect 29503 29121 29515 29155
rect 30650 29152 30656 29164
rect 30611 29124 30656 29152
rect 29457 29115 29515 29121
rect 24780 29056 25636 29084
rect 23845 29019 23903 29025
rect 23845 29016 23857 29019
rect 23400 28988 23857 29016
rect 19484 28920 22094 28948
rect 19484 28908 19490 28920
rect 22830 28908 22836 28960
rect 22888 28948 22894 28960
rect 23400 28948 23428 28988
rect 23845 28985 23857 28988
rect 23891 28985 23903 29019
rect 28368 29016 28396 29115
rect 30650 29112 30656 29124
rect 30708 29112 30714 29164
rect 30852 29161 30880 29192
rect 31481 29223 31539 29229
rect 31481 29189 31493 29223
rect 31527 29220 31539 29223
rect 32309 29223 32367 29229
rect 32309 29220 32321 29223
rect 31527 29192 32321 29220
rect 31527 29189 31539 29192
rect 31481 29183 31539 29189
rect 32309 29189 32321 29192
rect 32355 29189 32367 29223
rect 32309 29183 32367 29189
rect 33965 29223 34023 29229
rect 33965 29189 33977 29223
rect 34011 29220 34023 29223
rect 35802 29220 35808 29232
rect 34011 29192 35808 29220
rect 34011 29189 34023 29192
rect 33965 29183 34023 29189
rect 35802 29180 35808 29192
rect 35860 29180 35866 29232
rect 30837 29155 30895 29161
rect 30837 29121 30849 29155
rect 30883 29121 30895 29155
rect 30837 29115 30895 29121
rect 30929 29155 30987 29161
rect 30929 29121 30941 29155
rect 30975 29152 30987 29155
rect 31294 29152 31300 29164
rect 30975 29124 31300 29152
rect 30975 29121 30987 29124
rect 30929 29115 30987 29121
rect 31294 29112 31300 29124
rect 31352 29112 31358 29164
rect 31389 29153 31447 29159
rect 31389 29119 31401 29153
rect 31435 29119 31447 29153
rect 31389 29113 31447 29119
rect 29270 29084 29276 29096
rect 29231 29056 29276 29084
rect 29270 29044 29276 29056
rect 29328 29044 29334 29096
rect 31202 29044 31208 29096
rect 31260 29084 31266 29096
rect 31404 29084 31432 29113
rect 33778 29112 33784 29164
rect 33836 29152 33842 29164
rect 34422 29152 34428 29164
rect 33836 29124 34428 29152
rect 33836 29112 33842 29124
rect 34422 29112 34428 29124
rect 34480 29112 34486 29164
rect 34606 29152 34612 29164
rect 34567 29124 34612 29152
rect 34606 29112 34612 29124
rect 34664 29112 34670 29164
rect 35618 29112 35624 29164
rect 35676 29152 35682 29164
rect 35713 29155 35771 29161
rect 35713 29152 35725 29155
rect 35676 29124 35725 29152
rect 35676 29112 35682 29124
rect 35713 29121 35725 29124
rect 35759 29121 35771 29155
rect 37274 29152 37280 29164
rect 37235 29124 37280 29152
rect 35713 29115 35771 29121
rect 37274 29112 37280 29124
rect 37332 29112 37338 29164
rect 38105 29155 38163 29161
rect 38105 29121 38117 29155
rect 38151 29152 38163 29155
rect 38194 29152 38200 29164
rect 38151 29124 38200 29152
rect 38151 29121 38163 29124
rect 38105 29115 38163 29121
rect 38194 29112 38200 29124
rect 38252 29112 38258 29164
rect 31260 29056 31432 29084
rect 31260 29044 31266 29056
rect 31938 29044 31944 29096
rect 31996 29084 32002 29096
rect 32125 29087 32183 29093
rect 32125 29084 32137 29087
rect 31996 29056 32137 29084
rect 31996 29044 32002 29056
rect 32125 29053 32137 29056
rect 32171 29053 32183 29087
rect 32125 29047 32183 29053
rect 30374 29016 30380 29028
rect 28368 28988 30380 29016
rect 23845 28979 23903 28985
rect 30374 28976 30380 28988
rect 30432 29016 30438 29028
rect 30650 29016 30656 29028
rect 30432 28988 30656 29016
rect 30432 28976 30438 28988
rect 30650 28976 30656 28988
rect 30708 28976 30714 29028
rect 25130 28948 25136 28960
rect 22888 28920 23428 28948
rect 25091 28920 25136 28948
rect 22888 28908 22894 28920
rect 25130 28908 25136 28920
rect 25188 28908 25194 28960
rect 30926 28908 30932 28960
rect 30984 28948 30990 28960
rect 31846 28948 31852 28960
rect 30984 28920 31852 28948
rect 30984 28908 30990 28920
rect 31846 28908 31852 28920
rect 31904 28908 31910 28960
rect 34606 28948 34612 28960
rect 34567 28920 34612 28948
rect 34606 28908 34612 28920
rect 34664 28908 34670 28960
rect 35802 28948 35808 28960
rect 35763 28920 35808 28948
rect 35802 28908 35808 28920
rect 35860 28908 35866 28960
rect 36722 28948 36728 28960
rect 36683 28920 36728 28948
rect 36722 28908 36728 28920
rect 36780 28908 36786 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 1854 28704 1860 28756
rect 1912 28744 1918 28756
rect 2225 28747 2283 28753
rect 2225 28744 2237 28747
rect 1912 28716 2237 28744
rect 1912 28704 1918 28716
rect 2225 28713 2237 28716
rect 2271 28713 2283 28747
rect 2225 28707 2283 28713
rect 15930 28704 15936 28756
rect 15988 28744 15994 28756
rect 18049 28747 18107 28753
rect 15988 28716 18000 28744
rect 15988 28704 15994 28716
rect 17972 28676 18000 28716
rect 18049 28713 18061 28747
rect 18095 28744 18107 28747
rect 18230 28744 18236 28756
rect 18095 28716 18236 28744
rect 18095 28713 18107 28716
rect 18049 28707 18107 28713
rect 18230 28704 18236 28716
rect 18288 28704 18294 28756
rect 22649 28747 22707 28753
rect 22649 28713 22661 28747
rect 22695 28744 22707 28747
rect 22738 28744 22744 28756
rect 22695 28716 22744 28744
rect 22695 28713 22707 28716
rect 22649 28707 22707 28713
rect 22738 28704 22744 28716
rect 22796 28704 22802 28756
rect 24412 28716 25360 28744
rect 20438 28676 20444 28688
rect 17972 28648 20444 28676
rect 20438 28636 20444 28648
rect 20496 28676 20502 28688
rect 24412 28676 24440 28716
rect 20496 28648 24440 28676
rect 25332 28676 25360 28716
rect 25498 28704 25504 28756
rect 25556 28744 25562 28756
rect 25777 28747 25835 28753
rect 25777 28744 25789 28747
rect 25556 28716 25789 28744
rect 25556 28704 25562 28716
rect 25777 28713 25789 28716
rect 25823 28713 25835 28747
rect 27614 28744 27620 28756
rect 27575 28716 27620 28744
rect 25777 28707 25835 28713
rect 27614 28704 27620 28716
rect 27672 28704 27678 28756
rect 28258 28704 28264 28756
rect 28316 28744 28322 28756
rect 28537 28747 28595 28753
rect 28537 28744 28549 28747
rect 28316 28716 28549 28744
rect 28316 28704 28322 28716
rect 28537 28713 28549 28716
rect 28583 28713 28595 28747
rect 28537 28707 28595 28713
rect 28721 28747 28779 28753
rect 28721 28713 28733 28747
rect 28767 28744 28779 28747
rect 28902 28744 28908 28756
rect 28767 28716 28908 28744
rect 28767 28713 28779 28716
rect 28721 28707 28779 28713
rect 28902 28704 28908 28716
rect 28960 28704 28966 28756
rect 30926 28676 30932 28688
rect 25332 28648 30932 28676
rect 20496 28636 20502 28648
rect 30926 28636 30932 28648
rect 30984 28636 30990 28688
rect 31294 28636 31300 28688
rect 31352 28676 31358 28688
rect 31570 28676 31576 28688
rect 31352 28648 31576 28676
rect 31352 28636 31358 28648
rect 31570 28636 31576 28648
rect 31628 28676 31634 28688
rect 31628 28648 35664 28676
rect 31628 28636 31634 28648
rect 17313 28611 17371 28617
rect 17313 28577 17325 28611
rect 17359 28608 17371 28611
rect 18046 28608 18052 28620
rect 17359 28580 18052 28608
rect 17359 28577 17371 28580
rect 17313 28571 17371 28577
rect 18046 28568 18052 28580
rect 18104 28608 18110 28620
rect 19426 28608 19432 28620
rect 18104 28580 19432 28608
rect 18104 28568 18110 28580
rect 19426 28568 19432 28580
rect 19484 28568 19490 28620
rect 22462 28568 22468 28620
rect 22520 28608 22526 28620
rect 23474 28608 23480 28620
rect 22520 28580 23480 28608
rect 22520 28568 22526 28580
rect 23474 28568 23480 28580
rect 23532 28608 23538 28620
rect 24397 28611 24455 28617
rect 24397 28608 24409 28611
rect 23532 28580 24409 28608
rect 23532 28568 23538 28580
rect 24397 28577 24409 28580
rect 24443 28577 24455 28611
rect 32030 28608 32036 28620
rect 24397 28571 24455 28577
rect 26068 28580 32036 28608
rect 2314 28540 2320 28552
rect 2275 28512 2320 28540
rect 2314 28500 2320 28512
rect 2372 28500 2378 28552
rect 15286 28540 15292 28552
rect 15247 28512 15292 28540
rect 15286 28500 15292 28512
rect 15344 28500 15350 28552
rect 18138 28500 18144 28552
rect 18196 28540 18202 28552
rect 18279 28543 18337 28549
rect 18279 28540 18291 28543
rect 18196 28512 18291 28540
rect 18196 28500 18202 28512
rect 18279 28509 18291 28512
rect 18325 28509 18337 28543
rect 18279 28503 18337 28509
rect 18414 28543 18472 28549
rect 18414 28509 18426 28543
rect 18460 28509 18472 28543
rect 18414 28503 18472 28509
rect 4798 28432 4804 28484
rect 4856 28472 4862 28484
rect 9582 28472 9588 28484
rect 4856 28444 9588 28472
rect 4856 28432 4862 28444
rect 9582 28432 9588 28444
rect 9640 28432 9646 28484
rect 14642 28472 14648 28484
rect 14603 28444 14648 28472
rect 14642 28432 14648 28444
rect 14700 28432 14706 28484
rect 17068 28475 17126 28481
rect 17068 28441 17080 28475
rect 17114 28472 17126 28475
rect 17310 28472 17316 28484
rect 17114 28444 17316 28472
rect 17114 28441 17126 28444
rect 17068 28435 17126 28441
rect 17310 28432 17316 28444
rect 17368 28432 17374 28484
rect 18432 28472 18460 28503
rect 18506 28500 18512 28552
rect 18564 28549 18570 28552
rect 18564 28540 18572 28549
rect 18564 28512 18609 28540
rect 18564 28503 18572 28512
rect 18564 28500 18570 28503
rect 18690 28500 18696 28552
rect 18748 28540 18754 28552
rect 21450 28540 21456 28552
rect 18748 28512 21456 28540
rect 18748 28500 18754 28512
rect 21450 28500 21456 28512
rect 21508 28500 21514 28552
rect 22830 28500 22836 28552
rect 22888 28549 22894 28552
rect 22888 28543 22937 28549
rect 22888 28509 22891 28543
rect 22925 28509 22937 28543
rect 23014 28540 23020 28552
rect 22975 28512 23020 28540
rect 22888 28503 22937 28509
rect 22888 28500 22894 28503
rect 23014 28500 23020 28512
rect 23072 28500 23078 28552
rect 23106 28500 23112 28552
rect 23164 28540 23170 28552
rect 23164 28512 23209 28540
rect 23164 28500 23170 28512
rect 23290 28500 23296 28552
rect 23348 28540 23354 28552
rect 26068 28540 26096 28580
rect 32030 28568 32036 28580
rect 32088 28568 32094 28620
rect 33686 28608 33692 28620
rect 33647 28580 33692 28608
rect 33686 28568 33692 28580
rect 33744 28568 33750 28620
rect 34606 28608 34612 28620
rect 33796 28580 34612 28608
rect 33796 28552 33824 28580
rect 34606 28568 34612 28580
rect 34664 28608 34670 28620
rect 35636 28617 35664 28648
rect 35621 28611 35679 28617
rect 34664 28580 34744 28608
rect 34664 28568 34670 28580
rect 26878 28540 26884 28552
rect 23348 28512 26096 28540
rect 26839 28512 26884 28540
rect 23348 28500 23354 28512
rect 26878 28500 26884 28512
rect 26936 28500 26942 28552
rect 26973 28543 27031 28549
rect 26973 28509 26985 28543
rect 27019 28540 27031 28543
rect 27062 28540 27068 28552
rect 27019 28512 27068 28540
rect 27019 28509 27031 28512
rect 26973 28503 27031 28509
rect 27062 28500 27068 28512
rect 27120 28500 27126 28552
rect 27246 28500 27252 28552
rect 27304 28540 27310 28552
rect 27617 28543 27675 28549
rect 27617 28540 27629 28543
rect 27304 28512 27629 28540
rect 27304 28500 27310 28512
rect 27617 28509 27629 28512
rect 27663 28509 27675 28543
rect 27617 28503 27675 28509
rect 27801 28543 27859 28549
rect 27801 28509 27813 28543
rect 27847 28509 27859 28543
rect 33410 28540 33416 28552
rect 33371 28512 33416 28540
rect 27801 28503 27859 28509
rect 18782 28472 18788 28484
rect 18432 28444 18788 28472
rect 18782 28432 18788 28444
rect 18840 28432 18846 28484
rect 24664 28475 24722 28481
rect 24664 28441 24676 28475
rect 24710 28472 24722 28475
rect 24762 28472 24768 28484
rect 24710 28444 24768 28472
rect 24710 28441 24722 28444
rect 24664 28435 24722 28441
rect 24762 28432 24768 28444
rect 24820 28432 24826 28484
rect 27157 28475 27215 28481
rect 27157 28441 27169 28475
rect 27203 28472 27215 28475
rect 27816 28472 27844 28503
rect 33410 28500 33416 28512
rect 33468 28500 33474 28552
rect 33597 28543 33655 28549
rect 33597 28509 33609 28543
rect 33643 28509 33655 28543
rect 33778 28540 33784 28552
rect 33739 28512 33784 28540
rect 33597 28503 33655 28509
rect 28166 28472 28172 28484
rect 27203 28444 28172 28472
rect 27203 28441 27215 28444
rect 27157 28435 27215 28441
rect 28166 28432 28172 28444
rect 28224 28432 28230 28484
rect 28353 28475 28411 28481
rect 28353 28441 28365 28475
rect 28399 28472 28411 28475
rect 28442 28472 28448 28484
rect 28399 28444 28448 28472
rect 28399 28441 28411 28444
rect 28353 28435 28411 28441
rect 28442 28432 28448 28444
rect 28500 28472 28506 28484
rect 28810 28472 28816 28484
rect 28500 28444 28816 28472
rect 28500 28432 28506 28444
rect 28810 28432 28816 28444
rect 28868 28432 28874 28484
rect 33612 28472 33640 28503
rect 33778 28500 33784 28512
rect 33836 28500 33842 28552
rect 33962 28540 33968 28552
rect 33923 28512 33968 28540
rect 33962 28500 33968 28512
rect 34020 28500 34026 28552
rect 34716 28549 34744 28580
rect 35621 28577 35633 28611
rect 35667 28577 35679 28611
rect 35802 28608 35808 28620
rect 35763 28580 35808 28608
rect 35621 28571 35679 28577
rect 35802 28568 35808 28580
rect 35860 28568 35866 28620
rect 37090 28608 37096 28620
rect 37051 28580 37096 28608
rect 37090 28568 37096 28580
rect 37148 28568 37154 28620
rect 34701 28543 34759 28549
rect 34701 28509 34713 28543
rect 34747 28509 34759 28543
rect 34701 28503 34759 28509
rect 34790 28500 34796 28552
rect 34848 28540 34854 28552
rect 34977 28543 35035 28549
rect 34977 28540 34989 28543
rect 34848 28512 34989 28540
rect 34848 28500 34854 28512
rect 34977 28509 34989 28512
rect 35023 28509 35035 28543
rect 38102 28540 38108 28552
rect 38063 28512 38108 28540
rect 34977 28503 35035 28509
rect 38102 28500 38108 28512
rect 38160 28500 38166 28552
rect 34514 28472 34520 28484
rect 33612 28444 34520 28472
rect 34514 28432 34520 28444
rect 34572 28432 34578 28484
rect 15933 28407 15991 28413
rect 15933 28373 15945 28407
rect 15979 28404 15991 28407
rect 16666 28404 16672 28416
rect 15979 28376 16672 28404
rect 15979 28373 15991 28376
rect 15933 28367 15991 28373
rect 16666 28364 16672 28376
rect 16724 28404 16730 28416
rect 17586 28404 17592 28416
rect 16724 28376 17592 28404
rect 16724 28364 16730 28376
rect 17586 28364 17592 28376
rect 17644 28364 17650 28416
rect 28184 28404 28212 28432
rect 28553 28407 28611 28413
rect 28553 28404 28565 28407
rect 28184 28376 28565 28404
rect 28553 28373 28565 28376
rect 28599 28373 28611 28407
rect 28553 28367 28611 28373
rect 32858 28364 32864 28416
rect 32916 28404 32922 28416
rect 33229 28407 33287 28413
rect 33229 28404 33241 28407
rect 32916 28376 33241 28404
rect 32916 28364 32922 28376
rect 33229 28373 33241 28376
rect 33275 28373 33287 28407
rect 33229 28367 33287 28373
rect 33410 28364 33416 28416
rect 33468 28404 33474 28416
rect 34793 28407 34851 28413
rect 34793 28404 34805 28407
rect 33468 28376 34805 28404
rect 33468 28364 33474 28376
rect 34793 28373 34805 28376
rect 34839 28373 34851 28407
rect 34793 28367 34851 28373
rect 35161 28407 35219 28413
rect 35161 28373 35173 28407
rect 35207 28404 35219 28407
rect 36078 28404 36084 28416
rect 35207 28376 36084 28404
rect 35207 28373 35219 28376
rect 35161 28367 35219 28373
rect 36078 28364 36084 28376
rect 36136 28364 36142 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 17310 28200 17316 28212
rect 17271 28172 17316 28200
rect 17310 28160 17316 28172
rect 17368 28160 17374 28212
rect 22833 28203 22891 28209
rect 22833 28169 22845 28203
rect 22879 28200 22891 28203
rect 23106 28200 23112 28212
rect 22879 28172 23112 28200
rect 22879 28169 22891 28172
rect 22833 28163 22891 28169
rect 23106 28160 23112 28172
rect 23164 28160 23170 28212
rect 24762 28200 24768 28212
rect 24723 28172 24768 28200
rect 24762 28160 24768 28172
rect 24820 28160 24826 28212
rect 25225 28203 25283 28209
rect 25225 28169 25237 28203
rect 25271 28169 25283 28203
rect 27246 28200 27252 28212
rect 27207 28172 27252 28200
rect 25225 28163 25283 28169
rect 14182 28132 14188 28144
rect 12912 28104 14188 28132
rect 12912 28076 12940 28104
rect 14182 28092 14188 28104
rect 14240 28092 14246 28144
rect 19245 28135 19303 28141
rect 19245 28101 19257 28135
rect 19291 28132 19303 28135
rect 20254 28132 20260 28144
rect 19291 28104 20260 28132
rect 19291 28101 19303 28104
rect 19245 28095 19303 28101
rect 20254 28092 20260 28104
rect 20312 28132 20318 28144
rect 20622 28132 20628 28144
rect 20312 28104 20628 28132
rect 20312 28092 20318 28104
rect 20622 28092 20628 28104
rect 20680 28092 20686 28144
rect 21266 28092 21272 28144
rect 21324 28132 21330 28144
rect 21910 28132 21916 28144
rect 21324 28104 21916 28132
rect 21324 28092 21330 28104
rect 21910 28092 21916 28104
rect 21968 28132 21974 28144
rect 21968 28104 22048 28132
rect 21968 28092 21974 28104
rect 12894 28064 12900 28076
rect 12807 28036 12900 28064
rect 12894 28024 12900 28036
rect 12952 28024 12958 28076
rect 13633 28067 13691 28073
rect 13633 28064 13645 28067
rect 13096 28036 13645 28064
rect 13096 27937 13124 28036
rect 13633 28033 13645 28036
rect 13679 28064 13691 28067
rect 15197 28067 15255 28073
rect 15197 28064 15209 28067
rect 13679 28036 15209 28064
rect 13679 28033 13691 28036
rect 13633 28027 13691 28033
rect 15197 28033 15209 28036
rect 15243 28064 15255 28067
rect 15286 28064 15292 28076
rect 15243 28036 15292 28064
rect 15243 28033 15255 28036
rect 15197 28027 15255 28033
rect 15286 28024 15292 28036
rect 15344 28024 15350 28076
rect 17586 28064 17592 28076
rect 17547 28036 17592 28064
rect 17586 28024 17592 28036
rect 17644 28024 17650 28076
rect 17678 28067 17736 28073
rect 17678 28033 17690 28067
rect 17724 28033 17736 28067
rect 17678 28027 17736 28033
rect 14458 27996 14464 28008
rect 14419 27968 14464 27996
rect 14458 27956 14464 27968
rect 14516 27956 14522 28008
rect 15930 27996 15936 28008
rect 15891 27968 15936 27996
rect 15930 27956 15936 27968
rect 15988 27956 15994 28008
rect 17693 27940 17721 28027
rect 17770 28024 17776 28076
rect 17828 28073 17834 28076
rect 17828 28064 17836 28073
rect 17957 28067 18015 28073
rect 17828 28036 17873 28064
rect 17828 28027 17836 28036
rect 17957 28033 17969 28067
rect 18003 28064 18015 28067
rect 18690 28064 18696 28076
rect 18003 28036 18696 28064
rect 18003 28033 18015 28036
rect 17957 28027 18015 28033
rect 17828 28024 17834 28027
rect 18690 28024 18696 28036
rect 18748 28024 18754 28076
rect 19426 28024 19432 28076
rect 19484 28064 19490 28076
rect 20162 28073 20168 28076
rect 19889 28067 19947 28073
rect 19889 28064 19901 28067
rect 19484 28036 19901 28064
rect 19484 28024 19490 28036
rect 19889 28033 19901 28036
rect 19935 28033 19947 28067
rect 19889 28027 19947 28033
rect 20156 28027 20168 28073
rect 20220 28064 20226 28076
rect 20220 28036 20256 28064
rect 20162 28024 20168 28027
rect 20220 28024 20226 28036
rect 20898 28024 20904 28076
rect 20956 28064 20962 28076
rect 22020 28073 22048 28104
rect 21821 28067 21879 28073
rect 21821 28064 21833 28067
rect 20956 28036 21833 28064
rect 20956 28024 20962 28036
rect 21821 28033 21833 28036
rect 21867 28033 21879 28067
rect 21821 28027 21879 28033
rect 22005 28067 22063 28073
rect 22005 28033 22017 28067
rect 22051 28033 22063 28067
rect 22005 28027 22063 28033
rect 22278 28024 22284 28076
rect 22336 28064 22342 28076
rect 22649 28067 22707 28073
rect 22649 28064 22661 28067
rect 22336 28036 22661 28064
rect 22336 28024 22342 28036
rect 22649 28033 22661 28036
rect 22695 28033 22707 28067
rect 22649 28027 22707 28033
rect 22833 28067 22891 28073
rect 22833 28033 22845 28067
rect 22879 28033 22891 28067
rect 22833 28027 22891 28033
rect 24765 28067 24823 28073
rect 24765 28033 24777 28067
rect 24811 28064 24823 28067
rect 25240 28064 25268 28163
rect 27246 28160 27252 28172
rect 27304 28160 27310 28212
rect 28258 28200 28264 28212
rect 28219 28172 28264 28200
rect 28258 28160 28264 28172
rect 28316 28160 28322 28212
rect 31754 28160 31760 28212
rect 31812 28200 31818 28212
rect 32861 28203 32919 28209
rect 32861 28200 32873 28203
rect 31812 28172 32873 28200
rect 31812 28160 31818 28172
rect 32861 28169 32873 28172
rect 32907 28200 32919 28203
rect 33962 28200 33968 28212
rect 32907 28172 33968 28200
rect 32907 28169 32919 28172
rect 32861 28163 32919 28169
rect 33962 28160 33968 28172
rect 34020 28160 34026 28212
rect 25314 28092 25320 28144
rect 25372 28132 25378 28144
rect 25372 28101 25436 28132
rect 25372 28092 25375 28101
rect 24811 28036 25268 28064
rect 25363 28067 25375 28092
rect 25409 28070 25436 28101
rect 25498 28092 25504 28144
rect 25556 28132 25562 28144
rect 25593 28135 25651 28141
rect 25593 28132 25605 28135
rect 25556 28104 25605 28132
rect 25556 28092 25562 28104
rect 25593 28101 25605 28104
rect 25639 28101 25651 28135
rect 28442 28132 28448 28144
rect 28403 28104 28448 28132
rect 25593 28095 25651 28101
rect 28442 28092 28448 28104
rect 28500 28092 28506 28144
rect 38378 28132 38384 28144
rect 37292 28104 38384 28132
rect 25409 28067 25421 28070
rect 25363 28061 25421 28067
rect 24811 28033 24823 28036
rect 24765 28027 24823 28033
rect 22186 27956 22192 28008
rect 22244 27996 22250 28008
rect 22848 27996 22876 28027
rect 22244 27968 22876 27996
rect 22244 27956 22250 27968
rect 24302 27956 24308 28008
rect 24360 27996 24366 28008
rect 24489 27999 24547 28005
rect 24489 27996 24501 27999
rect 24360 27968 24501 27996
rect 24360 27956 24366 27968
rect 24489 27965 24501 27968
rect 24535 27965 24547 27999
rect 24489 27959 24547 27965
rect 24673 27999 24731 28005
rect 24673 27965 24685 27999
rect 24719 27996 24731 27999
rect 25130 27996 25136 28008
rect 24719 27968 25136 27996
rect 24719 27965 24731 27968
rect 24673 27959 24731 27965
rect 13081 27931 13139 27937
rect 13081 27897 13093 27931
rect 13127 27897 13139 27931
rect 13081 27891 13139 27897
rect 17678 27888 17684 27940
rect 17736 27888 17742 27940
rect 19426 27928 19432 27940
rect 19387 27900 19432 27928
rect 19426 27888 19432 27900
rect 19484 27888 19490 27940
rect 24504 27928 24532 27959
rect 25130 27956 25136 27968
rect 25188 27956 25194 28008
rect 25240 27996 25268 28036
rect 26878 28024 26884 28076
rect 26936 28064 26942 28076
rect 26973 28067 27031 28073
rect 26973 28064 26985 28067
rect 26936 28036 26985 28064
rect 26936 28024 26942 28036
rect 26973 28033 26985 28036
rect 27019 28033 27031 28067
rect 26973 28027 27031 28033
rect 27062 28024 27068 28076
rect 27120 28064 27126 28076
rect 28166 28064 28172 28076
rect 27120 28036 27165 28064
rect 28127 28036 28172 28064
rect 27120 28024 27126 28036
rect 28166 28024 28172 28036
rect 28224 28024 28230 28076
rect 28902 28064 28908 28076
rect 28863 28036 28908 28064
rect 28902 28024 28908 28036
rect 28960 28024 28966 28076
rect 30374 28024 30380 28076
rect 30432 28064 30438 28076
rect 31294 28064 31300 28076
rect 30432 28036 31300 28064
rect 30432 28024 30438 28036
rect 31294 28024 31300 28036
rect 31352 28024 31358 28076
rect 32950 28064 32956 28076
rect 32911 28036 32956 28064
rect 32950 28024 32956 28036
rect 33008 28024 33014 28076
rect 33410 28024 33416 28076
rect 33468 28064 33474 28076
rect 33505 28067 33563 28073
rect 33505 28064 33517 28067
rect 33468 28036 33517 28064
rect 33468 28024 33474 28036
rect 33505 28033 33517 28036
rect 33551 28033 33563 28067
rect 33778 28064 33784 28076
rect 33691 28036 33784 28064
rect 33505 28027 33563 28033
rect 33778 28024 33784 28036
rect 33836 28024 33842 28076
rect 33873 28067 33931 28073
rect 33873 28033 33885 28067
rect 33919 28064 33931 28067
rect 34514 28064 34520 28076
rect 33919 28036 34520 28064
rect 33919 28033 33931 28036
rect 33873 28027 33931 28033
rect 34514 28024 34520 28036
rect 34572 28024 34578 28076
rect 36722 28024 36728 28076
rect 36780 28064 36786 28076
rect 37292 28073 37320 28104
rect 38378 28092 38384 28104
rect 38436 28092 38442 28144
rect 37277 28067 37335 28073
rect 36780 28036 36825 28064
rect 36780 28024 36786 28036
rect 37277 28033 37289 28067
rect 37323 28033 37335 28067
rect 37277 28027 37335 28033
rect 37550 28024 37556 28076
rect 37608 28064 37614 28076
rect 37921 28067 37979 28073
rect 37921 28064 37933 28067
rect 37608 28036 37933 28064
rect 37608 28024 37614 28036
rect 37921 28033 37933 28036
rect 37967 28033 37979 28067
rect 37921 28027 37979 28033
rect 27080 27996 27108 28024
rect 25240 27968 27108 27996
rect 27154 27956 27160 28008
rect 27212 27996 27218 28008
rect 27249 27999 27307 28005
rect 27249 27996 27261 27999
rect 27212 27968 27261 27996
rect 27212 27956 27218 27968
rect 27249 27965 27261 27968
rect 27295 27965 27307 27999
rect 29181 27999 29239 28005
rect 29181 27996 29193 27999
rect 27249 27959 27307 27965
rect 27724 27968 29193 27996
rect 27724 27928 27752 27968
rect 29181 27965 29193 27968
rect 29227 27965 29239 27999
rect 29181 27959 29239 27965
rect 33597 27999 33655 28005
rect 33597 27965 33609 27999
rect 33643 27996 33655 27999
rect 33686 27996 33692 28008
rect 33643 27968 33692 27996
rect 33643 27965 33655 27968
rect 33597 27959 33655 27965
rect 24504 27900 27752 27928
rect 28445 27931 28503 27937
rect 28445 27897 28457 27931
rect 28491 27928 28503 27931
rect 28997 27931 29055 27937
rect 28997 27928 29009 27931
rect 28491 27900 29009 27928
rect 28491 27897 28503 27900
rect 28445 27891 28503 27897
rect 28997 27897 29009 27900
rect 29043 27897 29055 27931
rect 29196 27928 29224 27959
rect 33686 27956 33692 27968
rect 33744 27956 33750 28008
rect 31110 27928 31116 27940
rect 29196 27900 31116 27928
rect 28997 27891 29055 27897
rect 31110 27888 31116 27900
rect 31168 27928 31174 27940
rect 31481 27931 31539 27937
rect 31481 27928 31493 27931
rect 31168 27900 31493 27928
rect 31168 27888 31174 27900
rect 31481 27897 31493 27900
rect 31527 27897 31539 27931
rect 31481 27891 31539 27897
rect 33502 27888 33508 27940
rect 33560 27928 33566 27940
rect 33796 27928 33824 28024
rect 35710 27996 35716 28008
rect 35671 27968 35716 27996
rect 35710 27956 35716 27968
rect 35768 27956 35774 28008
rect 36541 27999 36599 28005
rect 36541 27965 36553 27999
rect 36587 27996 36599 27999
rect 38013 27999 38071 28005
rect 38013 27996 38025 27999
rect 36587 27968 38025 27996
rect 36587 27965 36599 27968
rect 36541 27959 36599 27965
rect 38013 27965 38025 27968
rect 38059 27965 38071 27999
rect 38013 27959 38071 27965
rect 33560 27900 33824 27928
rect 33560 27888 33566 27900
rect 21266 27860 21272 27872
rect 21227 27832 21272 27860
rect 21266 27820 21272 27832
rect 21324 27820 21330 27872
rect 22002 27860 22008 27872
rect 21963 27832 22008 27860
rect 22002 27820 22008 27832
rect 22060 27820 22066 27872
rect 25406 27860 25412 27872
rect 25367 27832 25412 27860
rect 25406 27820 25412 27832
rect 25464 27820 25470 27872
rect 29086 27860 29092 27872
rect 29047 27832 29092 27860
rect 29086 27820 29092 27832
rect 29144 27820 29150 27872
rect 34054 27860 34060 27872
rect 34015 27832 34060 27860
rect 34054 27820 34060 27832
rect 34112 27820 34118 27872
rect 37369 27863 37427 27869
rect 37369 27829 37381 27863
rect 37415 27860 37427 27863
rect 37918 27860 37924 27872
rect 37415 27832 37924 27860
rect 37415 27829 37427 27832
rect 37369 27823 37427 27829
rect 37918 27820 37924 27832
rect 37976 27820 37982 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 9582 27616 9588 27668
rect 9640 27656 9646 27668
rect 14642 27656 14648 27668
rect 9640 27628 14648 27656
rect 9640 27616 9646 27628
rect 14642 27616 14648 27628
rect 14700 27616 14706 27668
rect 17497 27659 17555 27665
rect 17497 27625 17509 27659
rect 17543 27656 17555 27659
rect 17770 27656 17776 27668
rect 17543 27628 17776 27656
rect 17543 27625 17555 27628
rect 17497 27619 17555 27625
rect 17770 27616 17776 27628
rect 17828 27616 17834 27668
rect 20162 27656 20168 27668
rect 20123 27628 20168 27656
rect 20162 27616 20168 27628
rect 20220 27616 20226 27668
rect 22186 27656 22192 27668
rect 20272 27628 22192 27656
rect 19426 27588 19432 27600
rect 18432 27560 19432 27588
rect 18432 27532 18460 27560
rect 19426 27548 19432 27560
rect 19484 27588 19490 27600
rect 20272 27588 20300 27628
rect 22186 27616 22192 27628
rect 22244 27616 22250 27668
rect 22278 27588 22284 27600
rect 19484 27560 20300 27588
rect 22239 27560 22284 27588
rect 19484 27548 19490 27560
rect 22278 27548 22284 27560
rect 22336 27548 22342 27600
rect 27338 27588 27344 27600
rect 27299 27560 27344 27588
rect 27338 27548 27344 27560
rect 27396 27548 27402 27600
rect 30834 27588 30840 27600
rect 27540 27560 30840 27588
rect 14826 27480 14832 27532
rect 14884 27520 14890 27532
rect 15105 27523 15163 27529
rect 15105 27520 15117 27523
rect 14884 27492 15117 27520
rect 14884 27480 14890 27492
rect 15105 27489 15117 27492
rect 15151 27520 15163 27523
rect 17494 27520 17500 27532
rect 15151 27492 17500 27520
rect 15151 27489 15163 27492
rect 15105 27483 15163 27489
rect 17494 27480 17500 27492
rect 17552 27480 17558 27532
rect 18414 27520 18420 27532
rect 17604 27492 18420 27520
rect 8021 27455 8079 27461
rect 8021 27421 8033 27455
rect 8067 27452 8079 27455
rect 8386 27452 8392 27464
rect 8067 27424 8392 27452
rect 8067 27421 8079 27424
rect 8021 27415 8079 27421
rect 8386 27412 8392 27424
rect 8444 27452 8450 27464
rect 12894 27452 12900 27464
rect 8444 27424 12900 27452
rect 8444 27412 8450 27424
rect 12894 27412 12900 27424
rect 12952 27412 12958 27464
rect 15286 27412 15292 27464
rect 15344 27452 15350 27464
rect 15473 27455 15531 27461
rect 15473 27452 15485 27455
rect 15344 27424 15485 27452
rect 15344 27412 15350 27424
rect 15473 27421 15485 27424
rect 15519 27452 15531 27455
rect 16209 27455 16267 27461
rect 16209 27452 16221 27455
rect 15519 27424 16221 27452
rect 15519 27421 15531 27424
rect 15473 27415 15531 27421
rect 16209 27421 16221 27424
rect 16255 27421 16267 27455
rect 16209 27415 16267 27421
rect 17218 27412 17224 27464
rect 17276 27452 17282 27464
rect 17604 27461 17632 27492
rect 18414 27480 18420 27492
rect 18472 27480 18478 27532
rect 19337 27523 19395 27529
rect 19337 27489 19349 27523
rect 19383 27520 19395 27523
rect 20070 27520 20076 27532
rect 19383 27492 20076 27520
rect 19383 27489 19395 27492
rect 19337 27483 19395 27489
rect 20070 27480 20076 27492
rect 20128 27480 20134 27532
rect 21266 27520 21272 27532
rect 20456 27492 21272 27520
rect 17405 27455 17463 27461
rect 17405 27452 17417 27455
rect 17276 27424 17417 27452
rect 17276 27412 17282 27424
rect 17405 27421 17417 27424
rect 17451 27421 17463 27455
rect 17405 27415 17463 27421
rect 17589 27455 17647 27461
rect 17589 27421 17601 27455
rect 17635 27421 17647 27455
rect 17589 27415 17647 27421
rect 18322 27412 18328 27464
rect 18380 27452 18386 27464
rect 19245 27455 19303 27461
rect 19245 27452 19257 27455
rect 18380 27424 19257 27452
rect 18380 27412 18386 27424
rect 19245 27421 19257 27424
rect 19291 27421 19303 27455
rect 19245 27415 19303 27421
rect 19429 27455 19487 27461
rect 19429 27421 19441 27455
rect 19475 27452 19487 27455
rect 19978 27452 19984 27464
rect 19475 27424 19984 27452
rect 19475 27421 19487 27424
rect 19429 27415 19487 27421
rect 19978 27412 19984 27424
rect 20036 27412 20042 27464
rect 20456 27461 20484 27492
rect 21266 27480 21272 27492
rect 21324 27480 21330 27532
rect 22002 27520 22008 27532
rect 21963 27492 22008 27520
rect 22002 27480 22008 27492
rect 22060 27480 22066 27532
rect 20441 27455 20499 27461
rect 20441 27421 20453 27455
rect 20487 27421 20499 27455
rect 20441 27415 20499 27421
rect 20533 27455 20591 27461
rect 20533 27421 20545 27455
rect 20579 27421 20591 27455
rect 20533 27415 20591 27421
rect 16758 27384 16764 27396
rect 16719 27356 16764 27384
rect 16758 27344 16764 27356
rect 16816 27344 16822 27396
rect 17770 27344 17776 27396
rect 17828 27384 17834 27396
rect 18782 27384 18788 27396
rect 17828 27356 18788 27384
rect 17828 27344 17834 27356
rect 18782 27344 18788 27356
rect 18840 27384 18846 27396
rect 20548 27384 20576 27415
rect 20622 27412 20628 27464
rect 20680 27452 20686 27464
rect 20809 27455 20867 27461
rect 20680 27424 20725 27452
rect 20680 27412 20686 27424
rect 20809 27421 20821 27455
rect 20855 27452 20867 27455
rect 21450 27452 21456 27464
rect 20855 27424 21456 27452
rect 20855 27421 20867 27424
rect 20809 27415 20867 27421
rect 21450 27412 21456 27424
rect 21508 27412 21514 27464
rect 21913 27455 21971 27461
rect 21913 27421 21925 27455
rect 21959 27452 21971 27455
rect 22094 27452 22100 27464
rect 21959 27424 22100 27452
rect 21959 27421 21971 27424
rect 21913 27415 21971 27421
rect 22094 27412 22100 27424
rect 22152 27412 22158 27464
rect 23198 27412 23204 27464
rect 23256 27452 23262 27464
rect 26142 27452 26148 27464
rect 23256 27424 26148 27452
rect 23256 27412 23262 27424
rect 26142 27412 26148 27424
rect 26200 27452 26206 27464
rect 27341 27455 27399 27461
rect 27341 27452 27353 27455
rect 26200 27424 27353 27452
rect 26200 27412 26206 27424
rect 27341 27421 27353 27424
rect 27387 27452 27399 27455
rect 27540 27452 27568 27560
rect 30834 27548 30840 27560
rect 30892 27548 30898 27600
rect 32677 27591 32735 27597
rect 32677 27557 32689 27591
rect 32723 27588 32735 27591
rect 32950 27588 32956 27600
rect 32723 27560 32956 27588
rect 32723 27557 32735 27560
rect 32677 27551 32735 27557
rect 32950 27548 32956 27560
rect 33008 27588 33014 27600
rect 33008 27560 33916 27588
rect 33008 27548 33014 27560
rect 28368 27492 31432 27520
rect 27387 27424 27568 27452
rect 27617 27455 27675 27461
rect 27387 27421 27399 27424
rect 27341 27415 27399 27421
rect 27617 27421 27629 27455
rect 27663 27452 27675 27455
rect 27706 27452 27712 27464
rect 27663 27424 27712 27452
rect 27663 27421 27675 27424
rect 27617 27415 27675 27421
rect 27706 27412 27712 27424
rect 27764 27452 27770 27464
rect 28166 27452 28172 27464
rect 27764 27424 28172 27452
rect 27764 27412 27770 27424
rect 28166 27412 28172 27424
rect 28224 27412 28230 27464
rect 23014 27384 23020 27396
rect 18840 27356 23020 27384
rect 18840 27344 18846 27356
rect 23014 27344 23020 27356
rect 23072 27344 23078 27396
rect 27525 27387 27583 27393
rect 27525 27353 27537 27387
rect 27571 27384 27583 27387
rect 27798 27384 27804 27396
rect 27571 27356 27804 27384
rect 27571 27353 27583 27356
rect 27525 27347 27583 27353
rect 27798 27344 27804 27356
rect 27856 27384 27862 27396
rect 28258 27384 28264 27396
rect 27856 27356 28264 27384
rect 27856 27344 27862 27356
rect 28258 27344 28264 27356
rect 28316 27344 28322 27396
rect 7834 27316 7840 27328
rect 7795 27288 7840 27316
rect 7834 27276 7840 27288
rect 7892 27276 7898 27328
rect 16776 27316 16804 27344
rect 28368 27316 28396 27492
rect 30653 27455 30711 27461
rect 30653 27421 30665 27455
rect 30699 27452 30711 27455
rect 30742 27452 30748 27464
rect 30699 27424 30748 27452
rect 30699 27421 30711 27424
rect 30653 27415 30711 27421
rect 30742 27412 30748 27424
rect 30800 27412 30806 27464
rect 31297 27455 31355 27461
rect 31297 27421 31309 27455
rect 31343 27421 31355 27455
rect 31404 27452 31432 27492
rect 33410 27480 33416 27532
rect 33468 27520 33474 27532
rect 33468 27492 33640 27520
rect 33468 27480 33474 27492
rect 33502 27452 33508 27464
rect 31404 27424 31754 27452
rect 33463 27424 33508 27452
rect 31297 27415 31355 27421
rect 31312 27384 31340 27415
rect 30760 27356 31340 27384
rect 16776 27288 28396 27316
rect 30650 27276 30656 27328
rect 30708 27316 30714 27328
rect 30760 27325 30788 27356
rect 31386 27344 31392 27396
rect 31444 27384 31450 27396
rect 31542 27387 31600 27393
rect 31542 27384 31554 27387
rect 31444 27356 31554 27384
rect 31444 27344 31450 27356
rect 31542 27353 31554 27356
rect 31588 27353 31600 27387
rect 31726 27384 31754 27424
rect 33502 27412 33508 27424
rect 33560 27412 33566 27464
rect 33612 27461 33640 27492
rect 33888 27461 33916 27560
rect 37182 27520 37188 27532
rect 37143 27492 37188 27520
rect 37182 27480 37188 27492
rect 37240 27480 37246 27532
rect 37918 27520 37924 27532
rect 37879 27492 37924 27520
rect 37918 27480 37924 27492
rect 37976 27480 37982 27532
rect 38102 27520 38108 27532
rect 38063 27492 38108 27520
rect 38102 27480 38108 27492
rect 38160 27480 38166 27532
rect 33597 27455 33655 27461
rect 33597 27421 33609 27455
rect 33643 27421 33655 27455
rect 33597 27415 33655 27421
rect 33781 27455 33839 27461
rect 33781 27421 33793 27455
rect 33827 27421 33839 27455
rect 33781 27415 33839 27421
rect 33873 27455 33931 27461
rect 33873 27421 33885 27455
rect 33919 27421 33931 27455
rect 33873 27415 33931 27421
rect 33796 27384 33824 27415
rect 34790 27384 34796 27396
rect 31726 27356 33732 27384
rect 33796 27356 34796 27384
rect 31542 27347 31600 27353
rect 30745 27319 30803 27325
rect 30745 27316 30757 27319
rect 30708 27288 30757 27316
rect 30708 27276 30714 27288
rect 30745 27285 30757 27288
rect 30791 27285 30803 27319
rect 33318 27316 33324 27328
rect 33279 27288 33324 27316
rect 30745 27279 30803 27285
rect 33318 27276 33324 27288
rect 33376 27276 33382 27328
rect 33704 27316 33732 27356
rect 34790 27344 34796 27356
rect 34848 27344 34854 27396
rect 37550 27316 37556 27328
rect 33704 27288 37556 27316
rect 37550 27276 37556 27288
rect 37608 27276 37614 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 8018 27072 8024 27124
rect 8076 27112 8082 27124
rect 17218 27112 17224 27124
rect 8076 27084 8432 27112
rect 17179 27084 17224 27112
rect 8076 27072 8082 27084
rect 8404 27053 8432 27084
rect 17218 27072 17224 27084
rect 17276 27072 17282 27124
rect 17770 27112 17776 27124
rect 17731 27084 17776 27112
rect 17770 27072 17776 27084
rect 17828 27072 17834 27124
rect 18506 27112 18512 27124
rect 18467 27084 18512 27112
rect 18506 27072 18512 27084
rect 18564 27072 18570 27124
rect 36265 27115 36323 27121
rect 18616 27084 36124 27112
rect 8389 27047 8447 27053
rect 8389 27013 8401 27047
rect 8435 27044 8447 27047
rect 18616 27044 18644 27084
rect 8435 27016 18644 27044
rect 19153 27047 19211 27053
rect 8435 27013 8447 27016
rect 8389 27007 8447 27013
rect 19153 27013 19165 27047
rect 19199 27044 19211 27047
rect 20254 27044 20260 27056
rect 19199 27016 20260 27044
rect 19199 27013 19211 27016
rect 19153 27007 19211 27013
rect 20254 27004 20260 27016
rect 20312 27004 20318 27056
rect 21085 27047 21143 27053
rect 21085 27013 21097 27047
rect 21131 27044 21143 27047
rect 22370 27044 22376 27056
rect 21131 27016 22376 27044
rect 21131 27013 21143 27016
rect 21085 27007 21143 27013
rect 22370 27004 22376 27016
rect 22428 27044 22434 27056
rect 26234 27044 26240 27056
rect 22428 27016 26240 27044
rect 22428 27004 22434 27016
rect 26234 27004 26240 27016
rect 26292 27004 26298 27056
rect 29086 27004 29092 27056
rect 29144 27044 29150 27056
rect 29558 27047 29616 27053
rect 29558 27044 29570 27047
rect 29144 27016 29570 27044
rect 29144 27004 29150 27016
rect 29558 27013 29570 27016
rect 29604 27013 29616 27047
rect 35710 27044 35716 27056
rect 29558 27007 29616 27013
rect 29656 27016 35716 27044
rect 7834 26936 7840 26988
rect 7892 26976 7898 26988
rect 8021 26979 8079 26985
rect 8021 26976 8033 26979
rect 7892 26948 8033 26976
rect 7892 26936 7898 26948
rect 8021 26945 8033 26948
rect 8067 26945 8079 26979
rect 14918 26976 14924 26988
rect 14879 26948 14924 26976
rect 8021 26939 8079 26945
rect 14918 26936 14924 26948
rect 14976 26936 14982 26988
rect 16850 26976 16856 26988
rect 16811 26948 16856 26976
rect 16850 26936 16856 26948
rect 16908 26936 16914 26988
rect 17865 26979 17923 26985
rect 17865 26945 17877 26979
rect 17911 26976 17923 26979
rect 18693 26979 18751 26985
rect 17911 26948 18368 26976
rect 17911 26945 17923 26948
rect 17865 26939 17923 26945
rect 15470 26908 15476 26920
rect 15431 26880 15476 26908
rect 15470 26868 15476 26880
rect 15528 26868 15534 26920
rect 16945 26911 17003 26917
rect 16945 26877 16957 26911
rect 16991 26908 17003 26911
rect 18046 26908 18052 26920
rect 16991 26880 18052 26908
rect 16991 26877 17003 26880
rect 16945 26871 17003 26877
rect 18046 26868 18052 26880
rect 18104 26868 18110 26920
rect 18340 26840 18368 26948
rect 18693 26945 18705 26979
rect 18739 26976 18751 26979
rect 20070 26976 20076 26988
rect 18739 26948 20076 26976
rect 18739 26945 18751 26948
rect 18693 26939 18751 26945
rect 20070 26936 20076 26948
rect 20128 26936 20134 26988
rect 21818 26976 21824 26988
rect 21779 26948 21824 26976
rect 21818 26936 21824 26948
rect 21876 26936 21882 26988
rect 21913 26979 21971 26985
rect 21913 26945 21925 26979
rect 21959 26945 21971 26979
rect 21913 26939 21971 26945
rect 18782 26868 18788 26920
rect 18840 26908 18846 26920
rect 21928 26908 21956 26939
rect 22002 26936 22008 26988
rect 22060 26976 22066 26988
rect 22097 26979 22155 26985
rect 22097 26976 22109 26979
rect 22060 26948 22109 26976
rect 22060 26936 22066 26948
rect 22097 26945 22109 26948
rect 22143 26945 22155 26979
rect 22097 26939 22155 26945
rect 22278 26936 22284 26988
rect 22336 26976 22342 26988
rect 22925 26979 22983 26985
rect 22925 26976 22937 26979
rect 22336 26948 22937 26976
rect 22336 26936 22342 26948
rect 22925 26945 22937 26948
rect 22971 26945 22983 26979
rect 22925 26939 22983 26945
rect 23017 26979 23075 26985
rect 23017 26945 23029 26979
rect 23063 26945 23075 26979
rect 23198 26976 23204 26988
rect 23159 26948 23204 26976
rect 23017 26939 23075 26945
rect 23032 26908 23060 26939
rect 23198 26936 23204 26948
rect 23256 26936 23262 26988
rect 25133 26979 25191 26985
rect 25133 26945 25145 26979
rect 25179 26945 25191 26979
rect 25406 26976 25412 26988
rect 25367 26948 25412 26976
rect 25133 26939 25191 26945
rect 23382 26908 23388 26920
rect 18840 26880 18885 26908
rect 21928 26880 23388 26908
rect 18840 26868 18846 26880
rect 22112 26852 22140 26880
rect 23382 26868 23388 26880
rect 23440 26868 23446 26920
rect 20162 26840 20168 26852
rect 18340 26812 20168 26840
rect 20162 26800 20168 26812
rect 20220 26840 20226 26852
rect 20441 26843 20499 26849
rect 20441 26840 20453 26843
rect 20220 26812 20453 26840
rect 20220 26800 20226 26812
rect 20441 26809 20453 26812
rect 20487 26809 20499 26843
rect 20441 26803 20499 26809
rect 22094 26800 22100 26852
rect 22152 26800 22158 26852
rect 25148 26840 25176 26939
rect 25406 26936 25412 26948
rect 25464 26936 25470 26988
rect 25866 26976 25872 26988
rect 25827 26948 25872 26976
rect 25866 26936 25872 26948
rect 25924 26936 25930 26988
rect 25961 26979 26019 26985
rect 25961 26945 25973 26979
rect 26007 26945 26019 26979
rect 26142 26976 26148 26988
rect 26103 26948 26148 26976
rect 25961 26939 26019 26945
rect 25424 26908 25452 26936
rect 25976 26908 26004 26939
rect 26142 26936 26148 26948
rect 26200 26936 26206 26988
rect 27338 26976 27344 26988
rect 27299 26948 27344 26976
rect 27338 26936 27344 26948
rect 27396 26936 27402 26988
rect 27525 26979 27583 26985
rect 27525 26945 27537 26979
rect 27571 26976 27583 26979
rect 27706 26976 27712 26988
rect 27571 26948 27712 26976
rect 27571 26945 27583 26948
rect 27525 26939 27583 26945
rect 27706 26936 27712 26948
rect 27764 26936 27770 26988
rect 29656 26976 29684 27016
rect 35710 27004 35716 27016
rect 35768 27004 35774 27056
rect 30374 26976 30380 26988
rect 27816 26948 29684 26976
rect 30335 26948 30380 26976
rect 26050 26908 26056 26920
rect 25424 26880 26056 26908
rect 26050 26868 26056 26880
rect 26108 26868 26114 26920
rect 27614 26908 27620 26920
rect 27575 26880 27620 26908
rect 27614 26868 27620 26880
rect 27672 26868 27678 26920
rect 26145 26843 26203 26849
rect 26145 26840 26157 26843
rect 25148 26812 26157 26840
rect 26145 26809 26157 26812
rect 26191 26809 26203 26843
rect 26145 26803 26203 26809
rect 26694 26800 26700 26852
rect 26752 26840 26758 26852
rect 27816 26840 27844 26948
rect 30374 26936 30380 26948
rect 30432 26936 30438 26988
rect 30558 26936 30564 26988
rect 30616 26976 30622 26988
rect 30834 26976 30840 26988
rect 30616 26948 30840 26976
rect 30616 26936 30622 26948
rect 30834 26936 30840 26948
rect 30892 26936 30898 26988
rect 34146 26936 34152 26988
rect 34204 26976 34210 26988
rect 35141 26979 35199 26985
rect 35141 26976 35153 26979
rect 34204 26948 35153 26976
rect 34204 26936 34210 26948
rect 35141 26945 35153 26948
rect 35187 26945 35199 26979
rect 36096 26976 36124 27084
rect 36265 27081 36277 27115
rect 36311 27081 36323 27115
rect 36265 27075 36323 27081
rect 36170 27004 36176 27056
rect 36228 27044 36234 27056
rect 36280 27044 36308 27075
rect 37829 27047 37887 27053
rect 37829 27044 37841 27047
rect 36228 27016 37841 27044
rect 36228 27004 36234 27016
rect 37829 27013 37841 27016
rect 37875 27013 37887 27047
rect 37829 27007 37887 27013
rect 37366 26976 37372 26988
rect 36096 26948 37372 26976
rect 35141 26939 35199 26945
rect 37366 26936 37372 26948
rect 37424 26936 37430 26988
rect 29822 26908 29828 26920
rect 29783 26880 29828 26908
rect 29822 26868 29828 26880
rect 29880 26908 29886 26920
rect 30650 26908 30656 26920
rect 29880 26880 30656 26908
rect 29880 26868 29886 26880
rect 30650 26868 30656 26880
rect 30708 26908 30714 26920
rect 30926 26908 30932 26920
rect 30708 26880 30932 26908
rect 30708 26868 30714 26880
rect 30926 26868 30932 26880
rect 30984 26908 30990 26920
rect 34885 26911 34943 26917
rect 34885 26908 34897 26911
rect 30984 26880 34897 26908
rect 30984 26868 30990 26880
rect 34885 26877 34897 26880
rect 34931 26877 34943 26911
rect 34885 26871 34943 26877
rect 37458 26868 37464 26920
rect 37516 26908 37522 26920
rect 37734 26908 37740 26920
rect 37516 26880 37740 26908
rect 37516 26868 37522 26880
rect 37734 26868 37740 26880
rect 37792 26868 37798 26920
rect 28442 26840 28448 26852
rect 26752 26812 27844 26840
rect 28403 26812 28448 26840
rect 26752 26800 26758 26812
rect 28442 26800 28448 26812
rect 28500 26800 28506 26852
rect 21174 26772 21180 26784
rect 21135 26744 21180 26772
rect 21174 26732 21180 26744
rect 21232 26732 21238 26784
rect 22002 26732 22008 26784
rect 22060 26772 22066 26784
rect 22281 26775 22339 26781
rect 22281 26772 22293 26775
rect 22060 26744 22293 26772
rect 22060 26732 22066 26744
rect 22281 26741 22293 26744
rect 22327 26741 22339 26775
rect 22281 26735 22339 26741
rect 22922 26732 22928 26784
rect 22980 26772 22986 26784
rect 23201 26775 23259 26781
rect 23201 26772 23213 26775
rect 22980 26744 23213 26772
rect 22980 26732 22986 26744
rect 23201 26741 23213 26744
rect 23247 26741 23259 26775
rect 24946 26772 24952 26784
rect 24907 26744 24952 26772
rect 23201 26735 23259 26741
rect 24946 26732 24952 26744
rect 25004 26732 25010 26784
rect 25314 26772 25320 26784
rect 25275 26744 25320 26772
rect 25314 26732 25320 26744
rect 25372 26772 25378 26784
rect 25866 26772 25872 26784
rect 25372 26744 25872 26772
rect 25372 26732 25378 26744
rect 25866 26732 25872 26744
rect 25924 26732 25930 26784
rect 27154 26772 27160 26784
rect 27115 26744 27160 26772
rect 27154 26732 27160 26744
rect 27212 26732 27218 26784
rect 32030 26732 32036 26784
rect 32088 26772 32094 26784
rect 32766 26772 32772 26784
rect 32088 26744 32772 26772
rect 32088 26732 32094 26744
rect 32766 26732 32772 26744
rect 32824 26772 32830 26784
rect 33502 26772 33508 26784
rect 32824 26744 33508 26772
rect 32824 26732 32830 26744
rect 33502 26732 33508 26744
rect 33560 26732 33566 26784
rect 34514 26732 34520 26784
rect 34572 26772 34578 26784
rect 35618 26772 35624 26784
rect 34572 26744 35624 26772
rect 34572 26732 34578 26744
rect 35618 26732 35624 26744
rect 35676 26772 35682 26784
rect 37737 26775 37795 26781
rect 37737 26772 37749 26775
rect 35676 26744 37749 26772
rect 35676 26732 35682 26744
rect 37737 26741 37749 26744
rect 37783 26741 37795 26775
rect 37737 26735 37795 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 15194 26528 15200 26580
rect 15252 26568 15258 26580
rect 15470 26568 15476 26580
rect 15252 26540 15476 26568
rect 15252 26528 15258 26540
rect 15470 26528 15476 26540
rect 15528 26568 15534 26580
rect 18693 26571 18751 26577
rect 15528 26540 17356 26568
rect 15528 26528 15534 26540
rect 16393 26503 16451 26509
rect 16393 26469 16405 26503
rect 16439 26500 16451 26503
rect 16850 26500 16856 26512
rect 16439 26472 16856 26500
rect 16439 26469 16451 26472
rect 16393 26463 16451 26469
rect 16850 26460 16856 26472
rect 16908 26500 16914 26512
rect 17328 26500 17356 26540
rect 18693 26537 18705 26571
rect 18739 26568 18751 26571
rect 18782 26568 18788 26580
rect 18739 26540 18788 26568
rect 18739 26537 18751 26540
rect 18693 26531 18751 26537
rect 18782 26528 18788 26540
rect 18840 26528 18846 26580
rect 18892 26540 20024 26568
rect 18892 26500 18920 26540
rect 16908 26472 17264 26500
rect 17328 26472 18920 26500
rect 19996 26500 20024 26540
rect 20622 26528 20628 26580
rect 20680 26568 20686 26580
rect 21085 26571 21143 26577
rect 21085 26568 21097 26571
rect 20680 26540 21097 26568
rect 20680 26528 20686 26540
rect 21085 26537 21097 26540
rect 21131 26537 21143 26571
rect 26050 26568 26056 26580
rect 21085 26531 21143 26537
rect 22066 26540 25636 26568
rect 26011 26540 26056 26568
rect 22066 26500 22094 26540
rect 19996 26472 22094 26500
rect 16908 26460 16914 26472
rect 16117 26435 16175 26441
rect 16117 26401 16129 26435
rect 16163 26432 16175 26435
rect 16574 26432 16580 26444
rect 16163 26404 16580 26432
rect 16163 26401 16175 26404
rect 16117 26395 16175 26401
rect 16574 26392 16580 26404
rect 16632 26392 16638 26444
rect 16025 26367 16083 26373
rect 16025 26333 16037 26367
rect 16071 26364 16083 26367
rect 16206 26364 16212 26376
rect 16071 26336 16212 26364
rect 16071 26333 16083 26336
rect 16025 26327 16083 26333
rect 16206 26324 16212 26336
rect 16264 26324 16270 26376
rect 17034 26364 17040 26376
rect 16995 26336 17040 26364
rect 17034 26324 17040 26336
rect 17092 26324 17098 26376
rect 17236 26373 17264 26472
rect 23382 26460 23388 26512
rect 23440 26500 23446 26512
rect 23753 26503 23811 26509
rect 23753 26500 23765 26503
rect 23440 26472 23765 26500
rect 23440 26460 23446 26472
rect 23753 26469 23765 26472
rect 23799 26469 23811 26503
rect 25608 26500 25636 26540
rect 26050 26528 26056 26540
rect 26108 26528 26114 26580
rect 27798 26528 27804 26580
rect 27856 26568 27862 26580
rect 28077 26571 28135 26577
rect 28077 26568 28089 26571
rect 27856 26540 28089 26568
rect 27856 26528 27862 26540
rect 28077 26537 28089 26540
rect 28123 26537 28135 26571
rect 31386 26568 31392 26580
rect 31347 26540 31392 26568
rect 28077 26531 28135 26537
rect 31386 26528 31392 26540
rect 31444 26528 31450 26580
rect 32950 26568 32956 26580
rect 31726 26540 32956 26568
rect 26694 26500 26700 26512
rect 25608 26472 26700 26500
rect 23753 26463 23811 26469
rect 26694 26460 26700 26472
rect 26752 26460 26758 26512
rect 30561 26503 30619 26509
rect 30561 26469 30573 26503
rect 30607 26500 30619 26503
rect 30650 26500 30656 26512
rect 30607 26472 30656 26500
rect 30607 26469 30619 26472
rect 30561 26463 30619 26469
rect 30650 26460 30656 26472
rect 30708 26460 30714 26512
rect 31726 26500 31754 26540
rect 32950 26528 32956 26540
rect 33008 26528 33014 26580
rect 34146 26568 34152 26580
rect 34107 26540 34152 26568
rect 34146 26528 34152 26540
rect 34204 26528 34210 26580
rect 30852 26472 31754 26500
rect 19334 26392 19340 26444
rect 19392 26432 19398 26444
rect 19521 26435 19579 26441
rect 19521 26432 19533 26435
rect 19392 26404 19533 26432
rect 19392 26392 19398 26404
rect 19521 26401 19533 26404
rect 19567 26401 19579 26435
rect 19521 26395 19579 26401
rect 19889 26435 19947 26441
rect 19889 26401 19901 26435
rect 19935 26432 19947 26435
rect 20070 26432 20076 26444
rect 19935 26404 20076 26432
rect 19935 26401 19947 26404
rect 19889 26395 19947 26401
rect 20070 26392 20076 26404
rect 20128 26392 20134 26444
rect 20254 26392 20260 26444
rect 20312 26432 20318 26444
rect 20441 26435 20499 26441
rect 20441 26432 20453 26435
rect 20312 26404 20453 26432
rect 20312 26392 20318 26404
rect 20441 26401 20453 26404
rect 20487 26401 20499 26435
rect 20441 26395 20499 26401
rect 20809 26435 20867 26441
rect 20809 26401 20821 26435
rect 20855 26432 20867 26435
rect 21545 26435 21603 26441
rect 21545 26432 21557 26435
rect 20855 26404 21557 26432
rect 20855 26401 20867 26404
rect 20809 26395 20867 26401
rect 21545 26401 21557 26404
rect 21591 26401 21603 26435
rect 21545 26395 21603 26401
rect 17221 26367 17279 26373
rect 17221 26333 17233 26367
rect 17267 26333 17279 26367
rect 17221 26327 17279 26333
rect 17313 26367 17371 26373
rect 17313 26333 17325 26367
rect 17359 26364 17371 26367
rect 18046 26364 18052 26376
rect 17359 26336 18052 26364
rect 17359 26333 17371 26336
rect 17313 26327 17371 26333
rect 18046 26324 18052 26336
rect 18104 26324 18110 26376
rect 18322 26364 18328 26376
rect 18283 26336 18328 26364
rect 18322 26324 18328 26336
rect 18380 26324 18386 26376
rect 19429 26367 19487 26373
rect 19429 26333 19441 26367
rect 19475 26364 19487 26367
rect 20901 26367 20959 26373
rect 19475 26336 20852 26364
rect 19475 26333 19487 26336
rect 19429 26327 19487 26333
rect 16850 26296 16856 26308
rect 16811 26268 16856 26296
rect 16850 26256 16856 26268
rect 16908 26256 16914 26308
rect 18506 26296 18512 26308
rect 18467 26268 18512 26296
rect 18506 26256 18512 26268
rect 18564 26256 18570 26308
rect 19242 26296 19248 26308
rect 19203 26268 19248 26296
rect 19242 26256 19248 26268
rect 19300 26256 19306 26308
rect 16942 26188 16948 26240
rect 17000 26228 17006 26240
rect 19444 26228 19472 26327
rect 20824 26308 20852 26336
rect 20901 26333 20913 26367
rect 20947 26364 20959 26367
rect 21082 26364 21088 26376
rect 20947 26336 21088 26364
rect 20947 26333 20959 26336
rect 20901 26327 20959 26333
rect 21082 26324 21088 26336
rect 21140 26324 21146 26376
rect 21174 26324 21180 26376
rect 21232 26364 21238 26376
rect 22373 26367 22431 26373
rect 22373 26364 22385 26367
rect 21232 26336 22385 26364
rect 21232 26324 21238 26336
rect 22373 26333 22385 26336
rect 22419 26364 22431 26367
rect 23474 26364 23480 26376
rect 22419 26336 23480 26364
rect 22419 26333 22431 26336
rect 22373 26327 22431 26333
rect 23474 26324 23480 26336
rect 23532 26364 23538 26376
rect 24394 26364 24400 26376
rect 23532 26336 24400 26364
rect 23532 26324 23538 26336
rect 24394 26324 24400 26336
rect 24452 26364 24458 26376
rect 24946 26373 24952 26376
rect 24673 26367 24731 26373
rect 24673 26364 24685 26367
rect 24452 26336 24685 26364
rect 24452 26324 24458 26336
rect 24673 26333 24685 26336
rect 24719 26333 24731 26367
rect 24940 26364 24952 26373
rect 24907 26336 24952 26364
rect 24673 26327 24731 26333
rect 24940 26327 24952 26336
rect 24946 26324 24952 26327
rect 25004 26324 25010 26376
rect 26697 26367 26755 26373
rect 26697 26333 26709 26367
rect 26743 26364 26755 26367
rect 29822 26364 29828 26376
rect 26743 26336 29828 26364
rect 26743 26333 26755 26336
rect 26697 26327 26755 26333
rect 29822 26324 29828 26336
rect 29880 26324 29886 26376
rect 30558 26364 30564 26376
rect 30519 26336 30564 26364
rect 30558 26324 30564 26336
rect 30616 26324 30622 26376
rect 30852 26373 30880 26472
rect 32122 26432 32128 26444
rect 31772 26404 32128 26432
rect 30837 26367 30895 26373
rect 30837 26333 30849 26367
rect 30883 26333 30895 26367
rect 31662 26364 31668 26376
rect 31623 26336 31668 26364
rect 30837 26327 30895 26333
rect 31662 26324 31668 26336
rect 31720 26324 31726 26376
rect 31772 26373 31800 26404
rect 32122 26392 32128 26404
rect 32180 26392 32186 26444
rect 33318 26432 33324 26444
rect 32600 26404 33324 26432
rect 31757 26367 31815 26373
rect 31757 26333 31769 26367
rect 31803 26333 31815 26367
rect 31757 26327 31815 26333
rect 31849 26367 31907 26373
rect 31849 26333 31861 26367
rect 31895 26333 31907 26367
rect 32030 26364 32036 26376
rect 31991 26336 32036 26364
rect 31849 26327 31907 26333
rect 20806 26256 20812 26308
rect 20864 26256 20870 26308
rect 21729 26299 21787 26305
rect 21729 26265 21741 26299
rect 21775 26265 21787 26299
rect 21729 26259 21787 26265
rect 17000 26200 19472 26228
rect 21744 26228 21772 26259
rect 21818 26256 21824 26308
rect 21876 26296 21882 26308
rect 21913 26299 21971 26305
rect 21913 26296 21925 26299
rect 21876 26268 21925 26296
rect 21876 26256 21882 26268
rect 21913 26265 21925 26268
rect 21959 26265 21971 26299
rect 21913 26259 21971 26265
rect 22640 26299 22698 26305
rect 22640 26265 22652 26299
rect 22686 26296 22698 26299
rect 22738 26296 22744 26308
rect 22686 26268 22744 26296
rect 22686 26265 22698 26268
rect 22640 26259 22698 26265
rect 22738 26256 22744 26268
rect 22796 26256 22802 26308
rect 26964 26299 27022 26305
rect 26964 26265 26976 26299
rect 27010 26296 27022 26299
rect 27154 26296 27160 26308
rect 27010 26268 27160 26296
rect 27010 26265 27022 26268
rect 26964 26259 27022 26265
rect 27154 26256 27160 26268
rect 27212 26256 27218 26308
rect 31864 26296 31892 26327
rect 32030 26324 32036 26336
rect 32088 26324 32094 26376
rect 32600 26373 32628 26404
rect 33318 26392 33324 26404
rect 33376 26392 33382 26444
rect 34514 26432 34520 26444
rect 33428 26404 33824 26432
rect 32585 26367 32643 26373
rect 32585 26333 32597 26367
rect 32631 26333 32643 26367
rect 32858 26364 32864 26376
rect 32819 26336 32864 26364
rect 32585 26327 32643 26333
rect 32858 26324 32864 26336
rect 32916 26324 32922 26376
rect 33042 26324 33048 26376
rect 33100 26364 33106 26376
rect 33428 26364 33456 26404
rect 33100 26336 33456 26364
rect 33100 26324 33106 26336
rect 33502 26324 33508 26376
rect 33560 26364 33566 26376
rect 33796 26373 33824 26404
rect 33888 26404 34520 26432
rect 33888 26373 33916 26404
rect 34514 26392 34520 26404
rect 34572 26392 34578 26444
rect 34698 26392 34704 26444
rect 34756 26432 34762 26444
rect 34885 26435 34943 26441
rect 34885 26432 34897 26435
rect 34756 26404 34897 26432
rect 34756 26392 34762 26404
rect 34885 26401 34897 26404
rect 34931 26401 34943 26435
rect 34885 26395 34943 26401
rect 35342 26392 35348 26444
rect 35400 26432 35406 26444
rect 35805 26435 35863 26441
rect 35805 26432 35817 26435
rect 35400 26404 35817 26432
rect 35400 26392 35406 26404
rect 35805 26401 35817 26404
rect 35851 26401 35863 26435
rect 36078 26432 36084 26444
rect 36039 26404 36084 26432
rect 35805 26395 35863 26401
rect 36078 26392 36084 26404
rect 36136 26392 36142 26444
rect 33689 26367 33747 26373
rect 33560 26336 33605 26364
rect 33560 26324 33566 26336
rect 33689 26333 33701 26367
rect 33735 26333 33747 26367
rect 33689 26327 33747 26333
rect 33781 26367 33839 26373
rect 33781 26333 33793 26367
rect 33827 26333 33839 26367
rect 33781 26327 33839 26333
rect 33873 26367 33931 26373
rect 33873 26333 33885 26367
rect 33919 26333 33931 26367
rect 33873 26327 33931 26333
rect 33226 26296 33232 26308
rect 31864 26268 33232 26296
rect 33226 26256 33232 26268
rect 33284 26256 33290 26308
rect 33704 26296 33732 26327
rect 34054 26324 34060 26376
rect 34112 26364 34118 26376
rect 34112 26336 34836 26364
rect 34112 26324 34118 26336
rect 34701 26299 34759 26305
rect 34701 26296 34713 26299
rect 33704 26268 34713 26296
rect 34701 26265 34713 26268
rect 34747 26265 34759 26299
rect 34808 26296 34836 26336
rect 34974 26324 34980 26376
rect 35032 26364 35038 26376
rect 36170 26364 36176 26376
rect 35032 26336 35077 26364
rect 36131 26336 36176 26364
rect 35032 26324 35038 26336
rect 36170 26324 36176 26336
rect 36228 26324 36234 26376
rect 37366 26364 37372 26376
rect 37327 26336 37372 26364
rect 37366 26324 37372 26336
rect 37424 26324 37430 26376
rect 35345 26299 35403 26305
rect 35345 26296 35357 26299
rect 34808 26268 35357 26296
rect 34701 26259 34759 26265
rect 35345 26265 35357 26268
rect 35391 26265 35403 26299
rect 37458 26296 37464 26308
rect 37419 26268 37464 26296
rect 35345 26259 35403 26265
rect 37458 26256 37464 26268
rect 37516 26256 37522 26308
rect 22002 26228 22008 26240
rect 21744 26200 22008 26228
rect 17000 26188 17006 26200
rect 22002 26188 22008 26200
rect 22060 26188 22066 26240
rect 30466 26188 30472 26240
rect 30524 26228 30530 26240
rect 30745 26231 30803 26237
rect 30745 26228 30757 26231
rect 30524 26200 30757 26228
rect 30524 26188 30530 26200
rect 30745 26197 30757 26200
rect 30791 26228 30803 26231
rect 31478 26228 31484 26240
rect 30791 26200 31484 26228
rect 30791 26197 30803 26200
rect 30745 26191 30803 26197
rect 31478 26188 31484 26200
rect 31536 26228 31542 26240
rect 32677 26231 32735 26237
rect 32677 26228 32689 26231
rect 31536 26200 32689 26228
rect 31536 26188 31542 26200
rect 32677 26197 32689 26200
rect 32723 26197 32735 26231
rect 32677 26191 32735 26197
rect 33045 26231 33103 26237
rect 33045 26197 33057 26231
rect 33091 26228 33103 26231
rect 34514 26228 34520 26240
rect 33091 26200 34520 26228
rect 33091 26197 33103 26200
rect 33045 26191 33103 26197
rect 34514 26188 34520 26200
rect 34572 26188 34578 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 17034 26024 17040 26036
rect 16995 25996 17040 26024
rect 17034 25984 17040 25996
rect 17092 25984 17098 26036
rect 18322 25984 18328 26036
rect 18380 26024 18386 26036
rect 18601 26027 18659 26033
rect 18601 26024 18613 26027
rect 18380 25996 18613 26024
rect 18380 25984 18386 25996
rect 18601 25993 18613 25996
rect 18647 25993 18659 26027
rect 18601 25987 18659 25993
rect 20809 26027 20867 26033
rect 20809 25993 20821 26027
rect 20855 26024 20867 26027
rect 20898 26024 20904 26036
rect 20855 25996 20904 26024
rect 20855 25993 20867 25996
rect 20809 25987 20867 25993
rect 20898 25984 20904 25996
rect 20956 25984 20962 26036
rect 21082 25984 21088 26036
rect 21140 26024 21146 26036
rect 21266 26024 21272 26036
rect 21140 25996 21272 26024
rect 21140 25984 21146 25996
rect 21266 25984 21272 25996
rect 21324 26024 21330 26036
rect 21913 26027 21971 26033
rect 21913 26024 21925 26027
rect 21324 25996 21925 26024
rect 21324 25984 21330 25996
rect 21913 25993 21925 25996
rect 21959 25993 21971 26027
rect 22738 26024 22744 26036
rect 22699 25996 22744 26024
rect 21913 25987 21971 25993
rect 22738 25984 22744 25996
rect 22796 25984 22802 26036
rect 26804 25996 31754 26024
rect 15838 25916 15844 25968
rect 15896 25956 15902 25968
rect 26804 25956 26832 25996
rect 15896 25928 26832 25956
rect 30316 25959 30374 25965
rect 15896 25916 15902 25928
rect 30316 25925 30328 25959
rect 30362 25956 30374 25959
rect 31021 25959 31079 25965
rect 31021 25956 31033 25959
rect 30362 25928 31033 25956
rect 30362 25925 30374 25928
rect 30316 25919 30374 25925
rect 31021 25925 31033 25928
rect 31067 25925 31079 25959
rect 31726 25956 31754 25996
rect 31846 25984 31852 26036
rect 31904 26024 31910 26036
rect 32122 26024 32128 26036
rect 31904 25996 32128 26024
rect 31904 25984 31910 25996
rect 32122 25984 32128 25996
rect 32180 26024 32186 26036
rect 33042 26024 33048 26036
rect 32180 25996 33048 26024
rect 32180 25984 32186 25996
rect 33042 25984 33048 25996
rect 33100 25984 33106 26036
rect 33226 26024 33232 26036
rect 33187 25996 33232 26024
rect 33226 25984 33232 25996
rect 33284 25984 33290 26036
rect 34333 26027 34391 26033
rect 34333 25993 34345 26027
rect 34379 26024 34391 26027
rect 34974 26024 34980 26036
rect 34379 25996 34980 26024
rect 34379 25993 34391 25996
rect 34333 25987 34391 25993
rect 34974 25984 34980 25996
rect 35032 25984 35038 26036
rect 31726 25928 37320 25956
rect 31021 25919 31079 25925
rect 16117 25891 16175 25897
rect 16117 25857 16129 25891
rect 16163 25888 16175 25891
rect 16666 25888 16672 25900
rect 16163 25860 16672 25888
rect 16163 25857 16175 25860
rect 16117 25851 16175 25857
rect 16666 25848 16672 25860
rect 16724 25848 16730 25900
rect 16853 25891 16911 25897
rect 16853 25857 16865 25891
rect 16899 25888 16911 25891
rect 16942 25888 16948 25900
rect 16899 25860 16948 25888
rect 16899 25857 16911 25860
rect 16853 25851 16911 25857
rect 16942 25848 16948 25860
rect 17000 25848 17006 25900
rect 18233 25891 18291 25897
rect 18233 25857 18245 25891
rect 18279 25888 18291 25891
rect 19150 25888 19156 25900
rect 18279 25860 19156 25888
rect 18279 25857 18291 25860
rect 18233 25851 18291 25857
rect 19150 25848 19156 25860
rect 19208 25848 19214 25900
rect 19245 25891 19303 25897
rect 19245 25857 19257 25891
rect 19291 25857 19303 25891
rect 19245 25851 19303 25857
rect 20717 25891 20775 25897
rect 20717 25857 20729 25891
rect 20763 25857 20775 25891
rect 20898 25888 20904 25900
rect 20859 25860 20904 25888
rect 20717 25851 20775 25857
rect 16574 25780 16580 25832
rect 16632 25820 16638 25832
rect 17862 25820 17868 25832
rect 16632 25792 17868 25820
rect 16632 25780 16638 25792
rect 17862 25780 17868 25792
rect 17920 25820 17926 25832
rect 18141 25823 18199 25829
rect 18141 25820 18153 25823
rect 17920 25792 18153 25820
rect 17920 25780 17926 25792
rect 18141 25789 18153 25792
rect 18187 25820 18199 25823
rect 19260 25820 19288 25851
rect 18187 25792 19288 25820
rect 18187 25789 18199 25792
rect 18141 25783 18199 25789
rect 19426 25780 19432 25832
rect 19484 25820 19490 25832
rect 19521 25823 19579 25829
rect 19521 25820 19533 25823
rect 19484 25792 19533 25820
rect 19484 25780 19490 25792
rect 19521 25789 19533 25792
rect 19567 25789 19579 25823
rect 19521 25783 19579 25789
rect 20732 25752 20760 25851
rect 20898 25848 20904 25860
rect 20956 25848 20962 25900
rect 21818 25888 21824 25900
rect 21731 25860 21824 25888
rect 21818 25848 21824 25860
rect 21876 25848 21882 25900
rect 22002 25888 22008 25900
rect 21963 25860 22008 25888
rect 22002 25848 22008 25860
rect 22060 25848 22066 25900
rect 22922 25888 22928 25900
rect 22883 25860 22928 25888
rect 22922 25848 22928 25860
rect 22980 25848 22986 25900
rect 23014 25848 23020 25900
rect 23072 25888 23078 25900
rect 23109 25891 23167 25897
rect 23109 25888 23121 25891
rect 23072 25860 23121 25888
rect 23072 25848 23078 25860
rect 23109 25857 23121 25860
rect 23155 25857 23167 25891
rect 25038 25888 25044 25900
rect 24999 25860 25044 25888
rect 23109 25851 23167 25857
rect 25038 25848 25044 25860
rect 25096 25848 25102 25900
rect 30650 25848 30656 25900
rect 30708 25888 30714 25900
rect 31205 25891 31263 25897
rect 31205 25888 31217 25891
rect 30708 25860 31217 25888
rect 30708 25848 30714 25860
rect 31205 25857 31217 25860
rect 31251 25857 31263 25891
rect 31205 25851 31263 25857
rect 31389 25891 31447 25897
rect 31389 25857 31401 25891
rect 31435 25888 31447 25891
rect 31846 25888 31852 25900
rect 31435 25860 31852 25888
rect 31435 25857 31447 25860
rect 31389 25851 31447 25857
rect 31846 25848 31852 25860
rect 31904 25848 31910 25900
rect 32309 25891 32367 25897
rect 32309 25888 32321 25891
rect 32048 25860 32321 25888
rect 20806 25780 20812 25832
rect 20864 25820 20870 25832
rect 21836 25820 21864 25848
rect 20864 25792 21864 25820
rect 23201 25823 23259 25829
rect 20864 25780 20870 25792
rect 23201 25789 23213 25823
rect 23247 25820 23259 25823
rect 23382 25820 23388 25832
rect 23247 25792 23388 25820
rect 23247 25789 23259 25792
rect 23201 25783 23259 25789
rect 23382 25780 23388 25792
rect 23440 25780 23446 25832
rect 25314 25820 25320 25832
rect 25275 25792 25320 25820
rect 25314 25780 25320 25792
rect 25372 25780 25378 25832
rect 30561 25823 30619 25829
rect 30561 25789 30573 25823
rect 30607 25820 30619 25823
rect 30926 25820 30932 25832
rect 30607 25792 30932 25820
rect 30607 25789 30619 25792
rect 30561 25783 30619 25789
rect 30926 25780 30932 25792
rect 30984 25780 30990 25832
rect 31478 25820 31484 25832
rect 31439 25792 31484 25820
rect 31478 25780 31484 25792
rect 31536 25820 31542 25832
rect 32048 25820 32076 25860
rect 32309 25857 32321 25860
rect 32355 25857 32367 25891
rect 33137 25891 33195 25897
rect 33137 25888 33149 25891
rect 32309 25851 32367 25857
rect 32692 25860 33149 25888
rect 32214 25820 32220 25832
rect 31536 25792 32076 25820
rect 32175 25792 32220 25820
rect 31536 25780 31542 25792
rect 32214 25780 32220 25792
rect 32272 25780 32278 25832
rect 22830 25752 22836 25764
rect 20732 25724 22836 25752
rect 22830 25712 22836 25724
rect 22888 25752 22894 25764
rect 23106 25752 23112 25764
rect 22888 25724 23112 25752
rect 22888 25712 22894 25724
rect 23106 25712 23112 25724
rect 23164 25712 23170 25764
rect 32692 25761 32720 25860
rect 33137 25857 33149 25860
rect 33183 25857 33195 25891
rect 33137 25851 33195 25857
rect 33321 25891 33379 25897
rect 33321 25857 33333 25891
rect 33367 25888 33379 25891
rect 33778 25888 33784 25900
rect 33367 25860 33784 25888
rect 33367 25857 33379 25860
rect 33321 25851 33379 25857
rect 33778 25848 33784 25860
rect 33836 25848 33842 25900
rect 34514 25888 34520 25900
rect 34475 25860 34520 25888
rect 34514 25848 34520 25860
rect 34572 25848 34578 25900
rect 34701 25891 34759 25897
rect 34701 25857 34713 25891
rect 34747 25888 34759 25891
rect 34790 25888 34796 25900
rect 34747 25860 34796 25888
rect 34747 25857 34759 25860
rect 34701 25851 34759 25857
rect 34790 25848 34796 25860
rect 34848 25888 34854 25900
rect 34974 25888 34980 25900
rect 34848 25860 34980 25888
rect 34848 25848 34854 25860
rect 34974 25848 34980 25860
rect 35032 25848 35038 25900
rect 35161 25891 35219 25897
rect 35161 25857 35173 25891
rect 35207 25857 35219 25891
rect 35342 25888 35348 25900
rect 35303 25860 35348 25888
rect 35161 25851 35219 25857
rect 34532 25820 34560 25848
rect 35176 25820 35204 25851
rect 35342 25848 35348 25860
rect 35400 25848 35406 25900
rect 37292 25897 37320 25928
rect 37277 25891 37335 25897
rect 37277 25857 37289 25891
rect 37323 25857 37335 25891
rect 37277 25851 37335 25857
rect 34532 25792 35204 25820
rect 32677 25755 32735 25761
rect 32677 25721 32689 25755
rect 32723 25721 32735 25755
rect 32677 25715 32735 25721
rect 16025 25687 16083 25693
rect 16025 25653 16037 25687
rect 16071 25684 16083 25687
rect 16206 25684 16212 25696
rect 16071 25656 16212 25684
rect 16071 25653 16083 25656
rect 16025 25647 16083 25653
rect 16206 25644 16212 25656
rect 16264 25644 16270 25696
rect 19058 25684 19064 25696
rect 19019 25656 19064 25684
rect 19058 25644 19064 25656
rect 19116 25644 19122 25696
rect 19334 25644 19340 25696
rect 19392 25684 19398 25696
rect 19429 25687 19487 25693
rect 19429 25684 19441 25687
rect 19392 25656 19441 25684
rect 19392 25644 19398 25656
rect 19429 25653 19441 25656
rect 19475 25653 19487 25687
rect 29178 25684 29184 25696
rect 29139 25656 29184 25684
rect 19429 25647 19487 25653
rect 29178 25644 29184 25656
rect 29236 25644 29242 25696
rect 34698 25644 34704 25696
rect 34756 25684 34762 25696
rect 35253 25687 35311 25693
rect 35253 25684 35265 25687
rect 34756 25656 35265 25684
rect 34756 25644 34762 25656
rect 35253 25653 35265 25656
rect 35299 25653 35311 25687
rect 36538 25684 36544 25696
rect 36499 25656 36544 25684
rect 35253 25647 35311 25653
rect 36538 25644 36544 25656
rect 36596 25644 36602 25696
rect 37369 25687 37427 25693
rect 37369 25653 37381 25687
rect 37415 25684 37427 25687
rect 37918 25684 37924 25696
rect 37415 25656 37924 25684
rect 37415 25653 37427 25656
rect 37369 25647 37427 25653
rect 37918 25644 37924 25656
rect 37976 25644 37982 25696
rect 38102 25684 38108 25696
rect 38063 25656 38108 25684
rect 38102 25644 38108 25656
rect 38160 25644 38166 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 18046 25480 18052 25492
rect 18007 25452 18052 25480
rect 18046 25440 18052 25452
rect 18104 25440 18110 25492
rect 18506 25440 18512 25492
rect 18564 25440 18570 25492
rect 25038 25440 25044 25492
rect 25096 25480 25102 25492
rect 25777 25483 25835 25489
rect 25777 25480 25789 25483
rect 25096 25452 25789 25480
rect 25096 25440 25102 25452
rect 25777 25449 25789 25452
rect 25823 25449 25835 25483
rect 32214 25480 32220 25492
rect 32175 25452 32220 25480
rect 25777 25443 25835 25449
rect 32214 25440 32220 25452
rect 32272 25440 32278 25492
rect 16761 25415 16819 25421
rect 16761 25381 16773 25415
rect 16807 25412 16819 25415
rect 16942 25412 16948 25424
rect 16807 25384 16948 25412
rect 16807 25381 16819 25384
rect 16761 25375 16819 25381
rect 16942 25372 16948 25384
rect 17000 25372 17006 25424
rect 18524 25412 18552 25440
rect 19978 25412 19984 25424
rect 18432 25384 19984 25412
rect 18322 25344 18328 25356
rect 18283 25316 18328 25344
rect 18322 25304 18328 25316
rect 18380 25304 18386 25356
rect 18432 25353 18460 25384
rect 19978 25372 19984 25384
rect 20036 25412 20042 25424
rect 20533 25415 20591 25421
rect 20533 25412 20545 25415
rect 20036 25384 20545 25412
rect 20036 25372 20042 25384
rect 20533 25381 20545 25384
rect 20579 25381 20591 25415
rect 20533 25375 20591 25381
rect 34514 25372 34520 25424
rect 34572 25412 34578 25424
rect 34572 25384 35112 25412
rect 34572 25372 34578 25384
rect 18417 25347 18475 25353
rect 18417 25313 18429 25347
rect 18463 25313 18475 25347
rect 18417 25307 18475 25313
rect 18509 25347 18567 25353
rect 18509 25313 18521 25347
rect 18555 25344 18567 25347
rect 19058 25344 19064 25356
rect 18555 25316 19064 25344
rect 18555 25313 18567 25316
rect 18509 25307 18567 25313
rect 19058 25304 19064 25316
rect 19116 25304 19122 25356
rect 20901 25347 20959 25353
rect 20901 25313 20913 25347
rect 20947 25344 20959 25347
rect 22002 25344 22008 25356
rect 20947 25316 22008 25344
rect 20947 25313 20959 25316
rect 20901 25307 20959 25313
rect 22002 25304 22008 25316
rect 22060 25304 22066 25356
rect 24394 25344 24400 25356
rect 24355 25316 24400 25344
rect 24394 25304 24400 25316
rect 24452 25304 24458 25356
rect 34790 25304 34796 25356
rect 34848 25344 34854 25356
rect 35084 25353 35112 25384
rect 34977 25347 35035 25353
rect 34977 25344 34989 25347
rect 34848 25316 34989 25344
rect 34848 25304 34854 25316
rect 34977 25313 34989 25316
rect 35023 25313 35035 25347
rect 34977 25307 35035 25313
rect 35069 25347 35127 25353
rect 35069 25313 35081 25347
rect 35115 25313 35127 25347
rect 37182 25344 37188 25356
rect 37143 25316 37188 25344
rect 35069 25307 35127 25313
rect 37182 25304 37188 25316
rect 37240 25304 37246 25356
rect 37918 25344 37924 25356
rect 37879 25316 37924 25344
rect 37918 25304 37924 25316
rect 37976 25304 37982 25356
rect 38102 25344 38108 25356
rect 38063 25316 38108 25344
rect 38102 25304 38108 25316
rect 38160 25304 38166 25356
rect 16574 25276 16580 25288
rect 16535 25248 16580 25276
rect 16574 25236 16580 25248
rect 16632 25236 16638 25288
rect 18230 25276 18236 25288
rect 18191 25248 18236 25276
rect 18230 25236 18236 25248
rect 18288 25236 18294 25288
rect 19334 25236 19340 25288
rect 19392 25276 19398 25288
rect 19429 25279 19487 25285
rect 19429 25276 19441 25279
rect 19392 25248 19441 25276
rect 19392 25236 19398 25248
rect 19429 25245 19441 25248
rect 19475 25245 19487 25279
rect 20714 25276 20720 25288
rect 20675 25248 20720 25276
rect 19429 25239 19487 25245
rect 20714 25236 20720 25248
rect 20772 25236 20778 25288
rect 20806 25236 20812 25288
rect 20864 25276 20870 25288
rect 20864 25248 20909 25276
rect 20864 25236 20870 25248
rect 20990 25236 20996 25288
rect 21048 25276 21054 25288
rect 21048 25248 21093 25276
rect 21048 25236 21054 25248
rect 29178 25236 29184 25288
rect 29236 25276 29242 25288
rect 29822 25276 29828 25288
rect 29236 25248 29828 25276
rect 29236 25236 29242 25248
rect 29822 25236 29828 25248
rect 29880 25276 29886 25288
rect 30377 25279 30435 25285
rect 30377 25276 30389 25279
rect 29880 25248 30389 25276
rect 29880 25236 29886 25248
rect 30377 25245 30389 25248
rect 30423 25245 30435 25279
rect 32030 25276 32036 25288
rect 31991 25248 32036 25276
rect 30377 25239 30435 25245
rect 32030 25236 32036 25248
rect 32088 25236 32094 25288
rect 32217 25279 32275 25285
rect 32217 25245 32229 25279
rect 32263 25276 32275 25279
rect 32858 25276 32864 25288
rect 32263 25248 32864 25276
rect 32263 25245 32275 25248
rect 32217 25239 32275 25245
rect 32858 25236 32864 25248
rect 32916 25236 32922 25288
rect 34882 25276 34888 25288
rect 34843 25248 34888 25276
rect 34882 25236 34888 25248
rect 34940 25236 34946 25288
rect 35161 25279 35219 25285
rect 35161 25245 35173 25279
rect 35207 25276 35219 25279
rect 35342 25276 35348 25288
rect 35207 25248 35348 25276
rect 35207 25245 35219 25248
rect 35161 25239 35219 25245
rect 35342 25236 35348 25248
rect 35400 25236 35406 25288
rect 24486 25168 24492 25220
rect 24544 25208 24550 25220
rect 24642 25211 24700 25217
rect 24642 25208 24654 25211
rect 24544 25180 24654 25208
rect 24544 25168 24550 25180
rect 24642 25177 24654 25180
rect 24688 25177 24700 25211
rect 24642 25171 24700 25177
rect 19150 25100 19156 25152
rect 19208 25140 19214 25152
rect 19337 25143 19395 25149
rect 19337 25140 19349 25143
rect 19208 25112 19349 25140
rect 19208 25100 19214 25112
rect 19337 25109 19349 25112
rect 19383 25109 19395 25143
rect 30466 25140 30472 25152
rect 30427 25112 30472 25140
rect 19337 25103 19395 25109
rect 30466 25100 30472 25112
rect 30524 25100 30530 25152
rect 34701 25143 34759 25149
rect 34701 25109 34713 25143
rect 34747 25140 34759 25143
rect 34790 25140 34796 25152
rect 34747 25112 34796 25140
rect 34747 25109 34759 25112
rect 34701 25103 34759 25109
rect 34790 25100 34796 25112
rect 34848 25100 34854 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 22021 24939 22079 24945
rect 22021 24936 22033 24939
rect 21008 24908 22033 24936
rect 15654 24800 15660 24812
rect 15615 24772 15660 24800
rect 15654 24760 15660 24772
rect 15712 24760 15718 24812
rect 15841 24803 15899 24809
rect 15841 24769 15853 24803
rect 15887 24800 15899 24803
rect 16850 24800 16856 24812
rect 15887 24772 16856 24800
rect 15887 24769 15899 24772
rect 15841 24763 15899 24769
rect 16850 24760 16856 24772
rect 16908 24760 16914 24812
rect 17862 24760 17868 24812
rect 17920 24800 17926 24812
rect 19705 24803 19763 24809
rect 19705 24800 19717 24803
rect 17920 24772 19717 24800
rect 17920 24760 17926 24772
rect 19705 24769 19717 24772
rect 19751 24769 19763 24803
rect 19705 24763 19763 24769
rect 19889 24803 19947 24809
rect 19889 24769 19901 24803
rect 19935 24769 19947 24803
rect 19889 24763 19947 24769
rect 19904 24732 19932 24763
rect 20714 24760 20720 24812
rect 20772 24800 20778 24812
rect 21008 24809 21036 24908
rect 22021 24905 22033 24908
rect 22067 24905 22079 24939
rect 24486 24936 24492 24948
rect 24447 24908 24492 24936
rect 22021 24899 22079 24905
rect 24486 24896 24492 24908
rect 24544 24896 24550 24948
rect 32030 24896 32036 24948
rect 32088 24936 32094 24948
rect 32217 24939 32275 24945
rect 32217 24936 32229 24939
rect 32088 24908 32229 24936
rect 32088 24896 32094 24908
rect 32217 24905 32229 24908
rect 32263 24905 32275 24939
rect 34777 24939 34835 24945
rect 34777 24936 34789 24939
rect 32217 24899 32275 24905
rect 34532 24908 34789 24936
rect 21821 24871 21879 24877
rect 21821 24868 21833 24871
rect 21192 24840 21833 24868
rect 20993 24803 21051 24809
rect 20993 24800 21005 24803
rect 20772 24772 21005 24800
rect 20772 24760 20778 24772
rect 20993 24769 21005 24772
rect 21039 24769 21051 24803
rect 20993 24763 21051 24769
rect 21082 24760 21088 24812
rect 21140 24800 21146 24812
rect 21192 24809 21220 24840
rect 21821 24837 21833 24840
rect 21867 24837 21879 24871
rect 34532 24868 34560 24908
rect 34777 24905 34789 24908
rect 34823 24936 34835 24939
rect 34882 24936 34888 24948
rect 34823 24908 34888 24936
rect 34823 24905 34835 24908
rect 34777 24899 34835 24905
rect 34882 24896 34888 24908
rect 34940 24936 34946 24948
rect 34940 24908 35572 24936
rect 34940 24896 34946 24908
rect 21821 24831 21879 24837
rect 27724 24840 28212 24868
rect 21177 24803 21235 24809
rect 21177 24800 21189 24803
rect 21140 24772 21189 24800
rect 21140 24760 21146 24772
rect 21177 24769 21189 24772
rect 21223 24769 21235 24803
rect 21177 24763 21235 24769
rect 21266 24760 21272 24812
rect 21324 24800 21330 24812
rect 24397 24803 24455 24809
rect 21324 24772 21369 24800
rect 21324 24760 21330 24772
rect 24397 24769 24409 24803
rect 24443 24769 24455 24803
rect 24397 24763 24455 24769
rect 24581 24803 24639 24809
rect 24581 24769 24593 24803
rect 24627 24800 24639 24803
rect 25314 24800 25320 24812
rect 24627 24772 25320 24800
rect 24627 24769 24639 24772
rect 24581 24763 24639 24769
rect 20530 24732 20536 24744
rect 19904 24704 20536 24732
rect 20530 24692 20536 24704
rect 20588 24732 20594 24744
rect 21634 24732 21640 24744
rect 20588 24704 21640 24732
rect 20588 24692 20594 24704
rect 21634 24692 21640 24704
rect 21692 24692 21698 24744
rect 24412 24732 24440 24763
rect 25314 24760 25320 24772
rect 25372 24760 25378 24812
rect 27338 24760 27344 24812
rect 27396 24800 27402 24812
rect 27724 24800 27752 24840
rect 27396 24772 27752 24800
rect 27801 24803 27859 24809
rect 27396 24760 27402 24772
rect 27801 24769 27813 24803
rect 27847 24769 27859 24803
rect 27801 24763 27859 24769
rect 27893 24803 27951 24809
rect 27893 24769 27905 24803
rect 27939 24769 27951 24803
rect 27893 24763 27951 24769
rect 25682 24732 25688 24744
rect 24412 24704 25688 24732
rect 25682 24692 25688 24704
rect 25740 24692 25746 24744
rect 27816 24664 27844 24763
rect 27908 24732 27936 24763
rect 27982 24760 27988 24812
rect 28040 24800 28046 24812
rect 28077 24803 28135 24809
rect 28077 24800 28089 24803
rect 28040 24772 28089 24800
rect 28040 24760 28046 24772
rect 28077 24769 28089 24772
rect 28123 24769 28135 24803
rect 28184 24800 28212 24840
rect 32048 24840 32260 24868
rect 28537 24803 28595 24809
rect 28537 24800 28549 24803
rect 28184 24772 28549 24800
rect 28077 24763 28135 24769
rect 28537 24769 28549 24772
rect 28583 24769 28595 24803
rect 28537 24763 28595 24769
rect 31754 24760 31760 24812
rect 31812 24800 31818 24812
rect 32048 24800 32076 24840
rect 31812 24772 32076 24800
rect 32125 24803 32183 24809
rect 31812 24760 31818 24772
rect 32125 24769 32137 24803
rect 32171 24769 32183 24803
rect 32232 24800 32260 24840
rect 33980 24840 34560 24868
rect 34977 24871 35035 24877
rect 32309 24803 32367 24809
rect 32309 24800 32321 24803
rect 32232 24772 32321 24800
rect 32125 24763 32183 24769
rect 32309 24769 32321 24772
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 28629 24735 28687 24741
rect 28629 24732 28641 24735
rect 27908 24704 28641 24732
rect 28629 24701 28641 24704
rect 28675 24732 28687 24735
rect 30006 24732 30012 24744
rect 28675 24704 30012 24732
rect 28675 24701 28687 24704
rect 28629 24695 28687 24701
rect 30006 24692 30012 24704
rect 30064 24692 30070 24744
rect 32140 24732 32168 24763
rect 32950 24760 32956 24812
rect 33008 24800 33014 24812
rect 33045 24803 33103 24809
rect 33045 24800 33057 24803
rect 33008 24772 33057 24800
rect 33008 24760 33014 24772
rect 33045 24769 33057 24772
rect 33091 24769 33103 24803
rect 33045 24763 33103 24769
rect 33229 24803 33287 24809
rect 33229 24769 33241 24803
rect 33275 24800 33287 24803
rect 33689 24803 33747 24809
rect 33689 24800 33701 24803
rect 33275 24772 33701 24800
rect 33275 24769 33287 24772
rect 33229 24763 33287 24769
rect 33689 24769 33701 24772
rect 33735 24769 33747 24803
rect 33689 24763 33747 24769
rect 33873 24803 33931 24809
rect 33873 24769 33885 24803
rect 33919 24800 33931 24803
rect 33980 24800 34008 24840
rect 34977 24837 34989 24871
rect 35023 24837 35035 24871
rect 34977 24831 35035 24837
rect 33919 24772 34008 24800
rect 34057 24803 34115 24809
rect 33919 24769 33931 24772
rect 33873 24763 33931 24769
rect 34057 24769 34069 24803
rect 34103 24769 34115 24803
rect 34057 24763 34115 24769
rect 33962 24732 33968 24744
rect 32140 24704 33968 24732
rect 33962 24692 33968 24704
rect 34020 24692 34026 24744
rect 34072 24732 34100 24763
rect 34146 24760 34152 24812
rect 34204 24800 34210 24812
rect 34992 24800 35020 24831
rect 34204 24772 34249 24800
rect 34532 24772 35020 24800
rect 34204 24760 34210 24772
rect 34532 24744 34560 24772
rect 34514 24732 34520 24744
rect 34072 24704 34520 24732
rect 34514 24692 34520 24704
rect 34572 24692 34578 24744
rect 35544 24741 35572 24908
rect 35894 24800 35900 24812
rect 35855 24772 35900 24800
rect 35894 24760 35900 24772
rect 35952 24760 35958 24812
rect 35529 24735 35587 24741
rect 35529 24701 35541 24735
rect 35575 24701 35587 24735
rect 35529 24695 35587 24701
rect 35989 24735 36047 24741
rect 35989 24701 36001 24735
rect 36035 24732 36047 24735
rect 36078 24732 36084 24744
rect 36035 24704 36084 24732
rect 36035 24701 36047 24704
rect 35989 24695 36047 24701
rect 36078 24692 36084 24704
rect 36136 24692 36142 24744
rect 29086 24664 29092 24676
rect 27816 24636 29092 24664
rect 29086 24624 29092 24636
rect 29144 24624 29150 24676
rect 33594 24624 33600 24676
rect 33652 24664 33658 24676
rect 34609 24667 34667 24673
rect 34609 24664 34621 24667
rect 33652 24636 34621 24664
rect 33652 24624 33658 24636
rect 34609 24633 34621 24636
rect 34655 24633 34667 24667
rect 34609 24627 34667 24633
rect 15749 24599 15807 24605
rect 15749 24565 15761 24599
rect 15795 24596 15807 24599
rect 15930 24596 15936 24608
rect 15795 24568 15936 24596
rect 15795 24565 15807 24568
rect 15749 24559 15807 24565
rect 15930 24556 15936 24568
rect 15988 24556 15994 24608
rect 20438 24556 20444 24608
rect 20496 24596 20502 24608
rect 20809 24599 20867 24605
rect 20809 24596 20821 24599
rect 20496 24568 20821 24596
rect 20496 24556 20502 24568
rect 20809 24565 20821 24568
rect 20855 24565 20867 24599
rect 20809 24559 20867 24565
rect 21266 24556 21272 24608
rect 21324 24596 21330 24608
rect 22005 24599 22063 24605
rect 22005 24596 22017 24599
rect 21324 24568 22017 24596
rect 21324 24556 21330 24568
rect 22005 24565 22017 24568
rect 22051 24565 22063 24599
rect 22186 24596 22192 24608
rect 22147 24568 22192 24596
rect 22005 24559 22063 24565
rect 22186 24556 22192 24568
rect 22244 24556 22250 24608
rect 28074 24596 28080 24608
rect 28035 24568 28080 24596
rect 28074 24556 28080 24568
rect 28132 24556 28138 24608
rect 29730 24556 29736 24608
rect 29788 24596 29794 24608
rect 30466 24596 30472 24608
rect 29788 24568 30472 24596
rect 29788 24556 29794 24568
rect 30466 24556 30472 24568
rect 30524 24556 30530 24608
rect 33137 24599 33195 24605
rect 33137 24565 33149 24599
rect 33183 24596 33195 24599
rect 33686 24596 33692 24608
rect 33183 24568 33692 24596
rect 33183 24565 33195 24568
rect 33137 24559 33195 24565
rect 33686 24556 33692 24568
rect 33744 24556 33750 24608
rect 34146 24556 34152 24608
rect 34204 24596 34210 24608
rect 34698 24596 34704 24608
rect 34204 24568 34704 24596
rect 34204 24556 34210 24568
rect 34698 24556 34704 24568
rect 34756 24596 34762 24608
rect 34793 24599 34851 24605
rect 34793 24596 34805 24599
rect 34756 24568 34805 24596
rect 34756 24556 34762 24568
rect 34793 24565 34805 24568
rect 34839 24565 34851 24599
rect 37826 24596 37832 24608
rect 37787 24568 37832 24596
rect 34793 24559 34851 24565
rect 37826 24556 37832 24568
rect 37884 24556 37890 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 15654 24352 15660 24404
rect 15712 24392 15718 24404
rect 15749 24395 15807 24401
rect 15749 24392 15761 24395
rect 15712 24364 15761 24392
rect 15712 24352 15718 24364
rect 15749 24361 15761 24364
rect 15795 24361 15807 24395
rect 15749 24355 15807 24361
rect 20901 24395 20959 24401
rect 20901 24361 20913 24395
rect 20947 24392 20959 24395
rect 20990 24392 20996 24404
rect 20947 24364 20996 24392
rect 20947 24361 20959 24364
rect 20901 24355 20959 24361
rect 15565 24259 15623 24265
rect 15565 24225 15577 24259
rect 15611 24225 15623 24259
rect 15565 24219 15623 24225
rect 15470 24188 15476 24200
rect 15431 24160 15476 24188
rect 15470 24148 15476 24160
rect 15528 24148 15534 24200
rect 15580 24120 15608 24219
rect 15764 24188 15792 24355
rect 20990 24352 20996 24364
rect 21048 24352 21054 24404
rect 21174 24352 21180 24404
rect 21232 24392 21238 24404
rect 21269 24395 21327 24401
rect 21269 24392 21281 24395
rect 21232 24364 21281 24392
rect 21232 24352 21238 24364
rect 21269 24361 21281 24364
rect 21315 24361 21327 24395
rect 33134 24392 33140 24404
rect 21269 24355 21327 24361
rect 21928 24364 33140 24392
rect 20349 24327 20407 24333
rect 20349 24293 20361 24327
rect 20395 24324 20407 24327
rect 20395 24296 21772 24324
rect 20395 24293 20407 24296
rect 20349 24287 20407 24293
rect 18325 24259 18383 24265
rect 18325 24225 18337 24259
rect 18371 24256 18383 24259
rect 19242 24256 19248 24268
rect 18371 24228 19248 24256
rect 18371 24225 18383 24228
rect 18325 24219 18383 24225
rect 19242 24216 19248 24228
rect 19300 24216 19306 24268
rect 21634 24256 21640 24268
rect 21100 24228 21640 24256
rect 16301 24191 16359 24197
rect 16301 24188 16313 24191
rect 15764 24160 16313 24188
rect 16301 24157 16313 24160
rect 16347 24157 16359 24191
rect 16301 24151 16359 24157
rect 16485 24191 16543 24197
rect 16485 24157 16497 24191
rect 16531 24188 16543 24191
rect 16850 24188 16856 24200
rect 16531 24160 16856 24188
rect 16531 24157 16543 24160
rect 16485 24151 16543 24157
rect 16850 24148 16856 24160
rect 16908 24148 16914 24200
rect 18230 24188 18236 24200
rect 18191 24160 18236 24188
rect 18230 24148 18236 24160
rect 18288 24148 18294 24200
rect 20162 24148 20168 24200
rect 20220 24188 20226 24200
rect 20257 24191 20315 24197
rect 20257 24188 20269 24191
rect 20220 24160 20269 24188
rect 20220 24148 20226 24160
rect 20257 24157 20269 24160
rect 20303 24157 20315 24191
rect 20438 24188 20444 24200
rect 20399 24160 20444 24188
rect 20257 24151 20315 24157
rect 20438 24148 20444 24160
rect 20496 24148 20502 24200
rect 21100 24197 21128 24228
rect 21634 24216 21640 24228
rect 21692 24216 21698 24268
rect 21085 24191 21143 24197
rect 21085 24157 21097 24191
rect 21131 24157 21143 24191
rect 21085 24151 21143 24157
rect 21361 24191 21419 24197
rect 21361 24157 21373 24191
rect 21407 24157 21419 24191
rect 21361 24151 21419 24157
rect 16942 24120 16948 24132
rect 15580 24092 16948 24120
rect 16942 24080 16948 24092
rect 17000 24080 17006 24132
rect 16022 24012 16028 24064
rect 16080 24052 16086 24064
rect 16669 24055 16727 24061
rect 16669 24052 16681 24055
rect 16080 24024 16681 24052
rect 16080 24012 16086 24024
rect 16669 24021 16681 24024
rect 16715 24021 16727 24055
rect 16669 24015 16727 24021
rect 18322 24012 18328 24064
rect 18380 24052 18386 24064
rect 18601 24055 18659 24061
rect 18601 24052 18613 24055
rect 18380 24024 18613 24052
rect 18380 24012 18386 24024
rect 18601 24021 18613 24024
rect 18647 24021 18659 24055
rect 21376 24052 21404 24151
rect 21744 24120 21772 24296
rect 21928 24197 21956 24364
rect 33134 24352 33140 24364
rect 33192 24392 33198 24404
rect 33410 24392 33416 24404
rect 33192 24364 33416 24392
rect 33192 24352 33198 24364
rect 33410 24352 33416 24364
rect 33468 24352 33474 24404
rect 35253 24395 35311 24401
rect 35253 24361 35265 24395
rect 35299 24392 35311 24395
rect 35342 24392 35348 24404
rect 35299 24364 35348 24392
rect 35299 24361 35311 24364
rect 35253 24355 35311 24361
rect 35342 24352 35348 24364
rect 35400 24352 35406 24404
rect 35618 24392 35624 24404
rect 35579 24364 35624 24392
rect 35618 24352 35624 24364
rect 35676 24352 35682 24404
rect 22186 24324 22192 24336
rect 22066 24296 22192 24324
rect 22066 24197 22094 24296
rect 22186 24284 22192 24296
rect 22244 24284 22250 24336
rect 25869 24327 25927 24333
rect 25869 24293 25881 24327
rect 25915 24324 25927 24327
rect 26605 24327 26663 24333
rect 26605 24324 26617 24327
rect 25915 24296 26617 24324
rect 25915 24293 25927 24296
rect 25869 24287 25927 24293
rect 26605 24293 26617 24296
rect 26651 24293 26663 24327
rect 27338 24324 27344 24336
rect 27299 24296 27344 24324
rect 26605 24287 26663 24293
rect 27338 24284 27344 24296
rect 27396 24284 27402 24336
rect 22278 24256 22284 24268
rect 22239 24228 22284 24256
rect 22278 24216 22284 24228
rect 22336 24216 22342 24268
rect 25682 24256 25688 24268
rect 25643 24228 25688 24256
rect 25682 24216 25688 24228
rect 25740 24216 25746 24268
rect 31754 24256 31760 24268
rect 29932 24228 31760 24256
rect 29932 24200 29960 24228
rect 31754 24216 31760 24228
rect 31812 24216 31818 24268
rect 33686 24256 33692 24268
rect 33647 24228 33692 24256
rect 33686 24216 33692 24228
rect 33744 24216 33750 24268
rect 33778 24216 33784 24268
rect 33836 24256 33842 24268
rect 36078 24256 36084 24268
rect 33836 24228 33881 24256
rect 35452 24228 36084 24256
rect 33836 24216 33842 24228
rect 35452 24200 35480 24228
rect 36078 24216 36084 24228
rect 36136 24216 36142 24268
rect 36265 24259 36323 24265
rect 36265 24225 36277 24259
rect 36311 24256 36323 24259
rect 36538 24256 36544 24268
rect 36311 24228 36544 24256
rect 36311 24225 36323 24228
rect 36265 24219 36323 24225
rect 36538 24216 36544 24228
rect 36596 24216 36602 24268
rect 38102 24256 38108 24268
rect 38063 24228 38108 24256
rect 38102 24216 38108 24228
rect 38160 24216 38166 24268
rect 21913 24191 21971 24197
rect 21913 24157 21925 24191
rect 21959 24157 21971 24191
rect 22066 24191 22127 24197
rect 22066 24160 22081 24191
rect 21913 24151 21971 24157
rect 22069 24157 22081 24160
rect 22115 24157 22127 24191
rect 22069 24151 22127 24157
rect 22189 24191 22247 24197
rect 22189 24157 22201 24191
rect 22235 24157 22247 24191
rect 22189 24151 22247 24157
rect 22465 24191 22523 24197
rect 22465 24157 22477 24191
rect 22511 24157 22523 24191
rect 22465 24151 22523 24157
rect 25961 24191 26019 24197
rect 25961 24157 25973 24191
rect 26007 24188 26019 24191
rect 26786 24188 26792 24200
rect 26007 24160 26792 24188
rect 26007 24157 26019 24160
rect 25961 24151 26019 24157
rect 22204 24120 22232 24151
rect 21744 24092 22232 24120
rect 22002 24052 22008 24064
rect 21376 24024 22008 24052
rect 18601 24015 18659 24021
rect 22002 24012 22008 24024
rect 22060 24052 22066 24064
rect 22480 24052 22508 24151
rect 26786 24148 26792 24160
rect 26844 24148 26850 24200
rect 26881 24191 26939 24197
rect 26881 24157 26893 24191
rect 26927 24188 26939 24191
rect 26970 24188 26976 24200
rect 26927 24160 26976 24188
rect 26927 24157 26939 24160
rect 26881 24151 26939 24157
rect 26970 24148 26976 24160
rect 27028 24148 27034 24200
rect 28074 24148 28080 24200
rect 28132 24188 28138 24200
rect 28454 24191 28512 24197
rect 28454 24188 28466 24191
rect 28132 24160 28466 24188
rect 28132 24148 28138 24160
rect 28454 24157 28466 24160
rect 28500 24157 28512 24191
rect 28454 24151 28512 24157
rect 28721 24191 28779 24197
rect 28721 24157 28733 24191
rect 28767 24157 28779 24191
rect 29546 24188 29552 24200
rect 29507 24160 29552 24188
rect 28721 24151 28779 24157
rect 26602 24120 26608 24132
rect 26563 24092 26608 24120
rect 26602 24080 26608 24092
rect 26660 24080 26666 24132
rect 28534 24080 28540 24132
rect 28592 24120 28598 24132
rect 28736 24120 28764 24151
rect 29546 24148 29552 24160
rect 29604 24148 29610 24200
rect 29730 24197 29736 24200
rect 29697 24191 29736 24197
rect 29697 24157 29709 24191
rect 29697 24151 29736 24157
rect 29730 24148 29736 24151
rect 29788 24148 29794 24200
rect 29914 24188 29920 24200
rect 29827 24160 29920 24188
rect 29914 24148 29920 24160
rect 29972 24148 29978 24200
rect 30006 24148 30012 24200
rect 30064 24197 30070 24200
rect 30064 24188 30072 24197
rect 30064 24160 30109 24188
rect 30064 24151 30072 24160
rect 30064 24148 30070 24151
rect 30742 24148 30748 24200
rect 30800 24188 30806 24200
rect 30837 24191 30895 24197
rect 30837 24188 30849 24191
rect 30800 24160 30849 24188
rect 30800 24148 30806 24160
rect 30837 24157 30849 24160
rect 30883 24157 30895 24191
rect 33410 24188 33416 24200
rect 33371 24160 33416 24188
rect 30837 24151 30895 24157
rect 33410 24148 33416 24160
rect 33468 24148 33474 24200
rect 33594 24188 33600 24200
rect 33555 24160 33600 24188
rect 33594 24148 33600 24160
rect 33652 24148 33658 24200
rect 33965 24191 34023 24197
rect 33965 24157 33977 24191
rect 34011 24157 34023 24191
rect 35434 24188 35440 24200
rect 35347 24160 35440 24188
rect 33965 24151 34023 24157
rect 28592 24092 28764 24120
rect 29825 24123 29883 24129
rect 28592 24080 28598 24092
rect 29825 24089 29837 24123
rect 29871 24120 29883 24123
rect 30098 24120 30104 24132
rect 29871 24092 30104 24120
rect 29871 24089 29883 24092
rect 29825 24083 29883 24089
rect 30098 24080 30104 24092
rect 30156 24080 30162 24132
rect 31018 24080 31024 24132
rect 31076 24120 31082 24132
rect 33980 24120 34008 24151
rect 35434 24148 35440 24160
rect 35492 24148 35498 24200
rect 35713 24191 35771 24197
rect 35713 24157 35725 24191
rect 35759 24188 35771 24191
rect 35894 24188 35900 24200
rect 35759 24160 35900 24188
rect 35759 24157 35771 24160
rect 35713 24151 35771 24157
rect 35728 24120 35756 24151
rect 35894 24148 35900 24160
rect 35952 24148 35958 24200
rect 31076 24092 35756 24120
rect 36449 24123 36507 24129
rect 31076 24080 31082 24092
rect 36449 24089 36461 24123
rect 36495 24120 36507 24123
rect 37458 24120 37464 24132
rect 36495 24092 37464 24120
rect 36495 24089 36507 24092
rect 36449 24083 36507 24089
rect 37458 24080 37464 24092
rect 37516 24080 37522 24132
rect 22646 24052 22652 24064
rect 22060 24024 22508 24052
rect 22607 24024 22652 24052
rect 22060 24012 22066 24024
rect 22646 24012 22652 24024
rect 22704 24012 22710 24064
rect 25958 24052 25964 24064
rect 25919 24024 25964 24052
rect 25958 24012 25964 24024
rect 26016 24012 26022 24064
rect 26789 24055 26847 24061
rect 26789 24021 26801 24055
rect 26835 24052 26847 24055
rect 27338 24052 27344 24064
rect 26835 24024 27344 24052
rect 26835 24021 26847 24024
rect 26789 24015 26847 24021
rect 27338 24012 27344 24024
rect 27396 24012 27402 24064
rect 30190 24052 30196 24064
rect 30151 24024 30196 24052
rect 30190 24012 30196 24024
rect 30248 24012 30254 24064
rect 30742 24052 30748 24064
rect 30703 24024 30748 24052
rect 30742 24012 30748 24024
rect 30800 24052 30806 24064
rect 32674 24052 32680 24064
rect 30800 24024 32680 24052
rect 30800 24012 30806 24024
rect 32674 24012 32680 24024
rect 32732 24012 32738 24064
rect 34149 24055 34207 24061
rect 34149 24021 34161 24055
rect 34195 24052 34207 24055
rect 35526 24052 35532 24064
rect 34195 24024 35532 24052
rect 34195 24021 34207 24024
rect 34149 24015 34207 24021
rect 35526 24012 35532 24024
rect 35584 24012 35590 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 15841 23851 15899 23857
rect 15841 23817 15853 23851
rect 15887 23817 15899 23851
rect 15841 23811 15899 23817
rect 15856 23780 15884 23811
rect 15930 23808 15936 23860
rect 15988 23848 15994 23860
rect 17681 23851 17739 23857
rect 15988 23820 16033 23848
rect 15988 23808 15994 23820
rect 17681 23817 17693 23851
rect 17727 23848 17739 23851
rect 18230 23848 18236 23860
rect 17727 23820 18236 23848
rect 17727 23817 17739 23820
rect 17681 23811 17739 23817
rect 18230 23808 18236 23820
rect 18288 23808 18294 23860
rect 18414 23848 18420 23860
rect 18375 23820 18420 23848
rect 18414 23808 18420 23820
rect 18472 23808 18478 23860
rect 21082 23848 21088 23860
rect 21043 23820 21088 23848
rect 21082 23808 21088 23820
rect 21140 23808 21146 23860
rect 22002 23808 22008 23860
rect 22060 23848 22066 23860
rect 22373 23851 22431 23857
rect 22373 23848 22385 23851
rect 22060 23820 22385 23848
rect 22060 23808 22066 23820
rect 22373 23817 22385 23820
rect 22419 23817 22431 23851
rect 22373 23811 22431 23817
rect 27338 23808 27344 23860
rect 27396 23848 27402 23860
rect 27709 23851 27767 23857
rect 27709 23848 27721 23851
rect 27396 23820 27721 23848
rect 27396 23808 27402 23820
rect 27709 23817 27721 23820
rect 27755 23817 27767 23851
rect 27709 23811 27767 23817
rect 27982 23808 27988 23860
rect 28040 23848 28046 23860
rect 28077 23851 28135 23857
rect 28077 23848 28089 23851
rect 28040 23820 28089 23848
rect 28040 23808 28046 23820
rect 28077 23817 28089 23820
rect 28123 23817 28135 23851
rect 28077 23811 28135 23817
rect 28534 23808 28540 23860
rect 28592 23848 28598 23860
rect 30742 23848 30748 23860
rect 28592 23820 30748 23848
rect 28592 23808 28598 23820
rect 30742 23808 30748 23820
rect 30800 23808 30806 23860
rect 34241 23851 34299 23857
rect 31726 23820 34192 23848
rect 16298 23780 16304 23792
rect 15856 23752 16304 23780
rect 16298 23740 16304 23752
rect 16356 23780 16362 23792
rect 18322 23780 18328 23792
rect 16356 23752 18184 23780
rect 18283 23752 18328 23780
rect 16356 23740 16362 23752
rect 15565 23715 15623 23721
rect 15565 23681 15577 23715
rect 15611 23712 15623 23715
rect 15838 23712 15844 23724
rect 15611 23684 15844 23712
rect 15611 23681 15623 23684
rect 15565 23675 15623 23681
rect 15838 23672 15844 23684
rect 15896 23672 15902 23724
rect 16022 23672 16028 23724
rect 16080 23712 16086 23724
rect 17313 23715 17371 23721
rect 16080 23684 16125 23712
rect 16080 23672 16086 23684
rect 17313 23681 17325 23715
rect 17359 23712 17371 23715
rect 17494 23712 17500 23724
rect 17359 23684 17500 23712
rect 17359 23681 17371 23684
rect 17313 23675 17371 23681
rect 17494 23672 17500 23684
rect 17552 23672 17558 23724
rect 18156 23712 18184 23752
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 20162 23780 20168 23792
rect 19260 23752 20168 23780
rect 19260 23721 19288 23752
rect 20162 23740 20168 23752
rect 20220 23740 20226 23792
rect 22646 23740 22652 23792
rect 22704 23780 22710 23792
rect 23486 23783 23544 23789
rect 23486 23780 23498 23783
rect 22704 23752 23498 23780
rect 22704 23740 22710 23752
rect 23486 23749 23498 23752
rect 23532 23749 23544 23783
rect 23486 23743 23544 23749
rect 25308 23783 25366 23789
rect 25308 23749 25320 23783
rect 25354 23780 25366 23783
rect 25958 23780 25964 23792
rect 25354 23752 25964 23780
rect 25354 23749 25366 23752
rect 25308 23743 25366 23749
rect 25958 23740 25964 23752
rect 26016 23740 26022 23792
rect 31726 23780 31754 23820
rect 29656 23752 31754 23780
rect 19245 23715 19303 23721
rect 19245 23712 19257 23715
rect 18156 23684 18368 23712
rect 17405 23647 17463 23653
rect 17405 23613 17417 23647
rect 17451 23644 17463 23647
rect 17862 23644 17868 23656
rect 17451 23616 17868 23644
rect 17451 23613 17463 23616
rect 17405 23607 17463 23613
rect 17862 23604 17868 23616
rect 17920 23604 17926 23656
rect 18340 23644 18368 23684
rect 18524 23684 19257 23712
rect 18524 23644 18552 23684
rect 19245 23681 19257 23684
rect 19291 23681 19303 23715
rect 19426 23712 19432 23724
rect 19387 23684 19432 23712
rect 19245 23675 19303 23681
rect 19426 23672 19432 23684
rect 19484 23672 19490 23724
rect 20898 23712 20904 23724
rect 20859 23684 20904 23712
rect 20898 23672 20904 23684
rect 20956 23672 20962 23724
rect 21085 23715 21143 23721
rect 21085 23681 21097 23715
rect 21131 23712 21143 23715
rect 21174 23712 21180 23724
rect 21131 23684 21180 23712
rect 21131 23681 21143 23684
rect 21085 23675 21143 23681
rect 21174 23672 21180 23684
rect 21232 23712 21238 23724
rect 22094 23712 22100 23724
rect 21232 23684 22100 23712
rect 21232 23672 21238 23684
rect 22094 23672 22100 23684
rect 22152 23672 22158 23724
rect 24302 23712 24308 23724
rect 22756 23684 24308 23712
rect 18340 23616 18552 23644
rect 18693 23647 18751 23653
rect 18693 23613 18705 23647
rect 18739 23644 18751 23647
rect 22756 23644 22784 23684
rect 24302 23672 24308 23684
rect 24360 23672 24366 23724
rect 26970 23712 26976 23724
rect 26931 23684 26976 23712
rect 26970 23672 26976 23684
rect 27028 23712 27034 23724
rect 27617 23715 27675 23721
rect 27617 23712 27629 23715
rect 27028 23684 27629 23712
rect 27028 23672 27034 23684
rect 27617 23681 27629 23684
rect 27663 23681 27675 23715
rect 27890 23712 27896 23724
rect 27851 23684 27896 23712
rect 27617 23675 27675 23681
rect 27890 23672 27896 23684
rect 27948 23672 27954 23724
rect 28537 23715 28595 23721
rect 28537 23681 28549 23715
rect 28583 23681 28595 23715
rect 28537 23675 28595 23681
rect 18739 23616 22784 23644
rect 23753 23647 23811 23653
rect 18739 23613 18751 23616
rect 18693 23607 18751 23613
rect 23753 23613 23765 23647
rect 23799 23644 23811 23647
rect 25038 23644 25044 23656
rect 23799 23616 25044 23644
rect 23799 23613 23811 23616
rect 23753 23607 23811 23613
rect 25038 23604 25044 23616
rect 25096 23604 25102 23656
rect 26602 23644 26608 23656
rect 26436 23616 26608 23644
rect 26436 23585 26464 23616
rect 26602 23604 26608 23616
rect 26660 23644 26666 23656
rect 27430 23644 27436 23656
rect 26660 23616 27436 23644
rect 26660 23604 26666 23616
rect 27430 23604 27436 23616
rect 27488 23644 27494 23656
rect 28552 23644 28580 23675
rect 28994 23672 29000 23724
rect 29052 23712 29058 23724
rect 29656 23721 29684 23752
rect 32306 23740 32312 23792
rect 32364 23780 32370 23792
rect 32585 23783 32643 23789
rect 32585 23780 32597 23783
rect 32364 23752 32597 23780
rect 32364 23740 32370 23752
rect 32585 23749 32597 23752
rect 32631 23780 32643 23783
rect 32950 23780 32956 23792
rect 32631 23752 32956 23780
rect 32631 23749 32643 23752
rect 32585 23743 32643 23749
rect 32950 23740 32956 23752
rect 33008 23780 33014 23792
rect 33413 23783 33471 23789
rect 33413 23780 33425 23783
rect 33008 23752 33425 23780
rect 33008 23740 33014 23752
rect 33413 23749 33425 23752
rect 33459 23749 33471 23783
rect 33413 23743 33471 23749
rect 34164 23780 34192 23820
rect 34241 23817 34253 23851
rect 34287 23848 34299 23851
rect 34514 23848 34520 23860
rect 34287 23820 34520 23848
rect 34287 23817 34299 23820
rect 34241 23811 34299 23817
rect 34514 23808 34520 23820
rect 34572 23808 34578 23860
rect 35618 23848 35624 23860
rect 34624 23820 35624 23848
rect 34624 23780 34652 23820
rect 35618 23808 35624 23820
rect 35676 23808 35682 23860
rect 35894 23808 35900 23860
rect 35952 23848 35958 23860
rect 36633 23851 36691 23857
rect 36633 23848 36645 23851
rect 35952 23820 36645 23848
rect 35952 23808 35958 23820
rect 36633 23817 36645 23820
rect 36679 23817 36691 23851
rect 36633 23811 36691 23817
rect 35526 23789 35532 23792
rect 35520 23780 35532 23789
rect 34164 23752 34652 23780
rect 35487 23752 35532 23780
rect 29641 23715 29699 23721
rect 29641 23712 29653 23715
rect 29052 23684 29653 23712
rect 29052 23672 29058 23684
rect 29641 23681 29653 23684
rect 29687 23681 29699 23715
rect 29914 23712 29920 23724
rect 29875 23684 29920 23712
rect 29641 23675 29699 23681
rect 29914 23672 29920 23684
rect 29972 23672 29978 23724
rect 30006 23672 30012 23724
rect 30064 23712 30070 23724
rect 30190 23712 30196 23724
rect 30064 23684 30109 23712
rect 30151 23684 30196 23712
rect 30064 23672 30070 23684
rect 30190 23672 30196 23684
rect 30248 23672 30254 23724
rect 33594 23712 33600 23724
rect 33507 23684 33600 23712
rect 33594 23672 33600 23684
rect 33652 23712 33658 23724
rect 34054 23712 34060 23724
rect 33652 23684 34060 23712
rect 33652 23672 33658 23684
rect 34054 23672 34060 23684
rect 34112 23672 34118 23724
rect 34164 23721 34192 23752
rect 35520 23743 35532 23752
rect 35526 23740 35532 23743
rect 35584 23740 35590 23792
rect 34149 23715 34207 23721
rect 34333 23718 34391 23721
rect 34149 23681 34161 23715
rect 34195 23681 34207 23715
rect 34149 23675 34207 23681
rect 34256 23715 34391 23718
rect 34256 23690 34345 23715
rect 27488 23616 28580 23644
rect 28629 23647 28687 23653
rect 27488 23604 27494 23616
rect 28629 23613 28641 23647
rect 28675 23644 28687 23647
rect 28810 23644 28816 23656
rect 28675 23616 28816 23644
rect 28675 23613 28687 23616
rect 28629 23607 28687 23613
rect 28810 23604 28816 23616
rect 28868 23644 28874 23656
rect 29825 23647 29883 23653
rect 29825 23644 29837 23647
rect 28868 23616 29837 23644
rect 28868 23604 28874 23616
rect 29825 23613 29837 23616
rect 29871 23613 29883 23647
rect 29825 23607 29883 23613
rect 33962 23604 33968 23656
rect 34020 23644 34026 23656
rect 34256 23644 34284 23690
rect 34333 23681 34345 23690
rect 34379 23681 34391 23715
rect 34333 23675 34391 23681
rect 35253 23715 35311 23721
rect 35253 23681 35265 23715
rect 35299 23712 35311 23715
rect 35342 23712 35348 23724
rect 35299 23684 35348 23712
rect 35299 23681 35311 23684
rect 35253 23675 35311 23681
rect 34020 23616 34284 23644
rect 34020 23604 34026 23616
rect 18601 23579 18659 23585
rect 18601 23545 18613 23579
rect 18647 23576 18659 23579
rect 19245 23579 19303 23585
rect 19245 23576 19257 23579
rect 18647 23548 19257 23576
rect 18647 23545 18659 23548
rect 18601 23539 18659 23545
rect 19245 23545 19257 23548
rect 19291 23545 19303 23579
rect 19245 23539 19303 23545
rect 26421 23579 26479 23585
rect 26421 23545 26433 23579
rect 26467 23545 26479 23579
rect 26421 23539 26479 23545
rect 27065 23579 27123 23585
rect 27065 23545 27077 23579
rect 27111 23576 27123 23579
rect 29086 23576 29092 23588
rect 27111 23548 29092 23576
rect 27111 23545 27123 23548
rect 27065 23539 27123 23545
rect 29086 23536 29092 23548
rect 29144 23576 29150 23588
rect 30098 23576 30104 23588
rect 29144 23548 30104 23576
rect 29144 23536 29150 23548
rect 30098 23536 30104 23548
rect 30156 23536 30162 23588
rect 32769 23579 32827 23585
rect 32769 23545 32781 23579
rect 32815 23576 32827 23579
rect 32858 23576 32864 23588
rect 32815 23548 32864 23576
rect 32815 23545 32827 23548
rect 32769 23539 32827 23545
rect 32858 23536 32864 23548
rect 32916 23536 32922 23588
rect 15562 23508 15568 23520
rect 15523 23480 15568 23508
rect 15562 23468 15568 23480
rect 15620 23468 15626 23520
rect 15654 23468 15660 23520
rect 15712 23508 15718 23520
rect 18690 23508 18696 23520
rect 15712 23480 15757 23508
rect 18651 23480 18696 23508
rect 15712 23468 15718 23480
rect 18690 23468 18696 23480
rect 18748 23468 18754 23520
rect 29457 23511 29515 23517
rect 29457 23477 29469 23511
rect 29503 23508 29515 23511
rect 29638 23508 29644 23520
rect 29503 23480 29644 23508
rect 29503 23477 29515 23480
rect 29457 23471 29515 23477
rect 29638 23468 29644 23480
rect 29696 23468 29702 23520
rect 32674 23468 32680 23520
rect 32732 23508 32738 23520
rect 35268 23508 35296 23675
rect 35342 23672 35348 23684
rect 35400 23672 35406 23724
rect 37274 23672 37280 23724
rect 37332 23712 37338 23724
rect 37369 23715 37427 23721
rect 37369 23712 37381 23715
rect 37332 23684 37381 23712
rect 37332 23672 37338 23684
rect 37369 23681 37381 23684
rect 37415 23712 37427 23715
rect 38286 23712 38292 23724
rect 37415 23684 38292 23712
rect 37415 23681 37427 23684
rect 37369 23675 37427 23681
rect 38286 23672 38292 23684
rect 38344 23672 38350 23724
rect 32732 23480 35296 23508
rect 37461 23511 37519 23517
rect 32732 23468 32738 23480
rect 37461 23477 37473 23511
rect 37507 23508 37519 23511
rect 37918 23508 37924 23520
rect 37507 23480 37924 23508
rect 37507 23477 37519 23480
rect 37461 23471 37519 23477
rect 37918 23468 37924 23480
rect 37976 23468 37982 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 15654 23264 15660 23316
rect 15712 23304 15718 23316
rect 16301 23307 16359 23313
rect 16301 23304 16313 23307
rect 15712 23276 16313 23304
rect 15712 23264 15718 23276
rect 16301 23273 16313 23276
rect 16347 23273 16359 23307
rect 16301 23267 16359 23273
rect 17494 23264 17500 23316
rect 17552 23304 17558 23316
rect 19337 23307 19395 23313
rect 19337 23304 19349 23307
rect 17552 23276 19349 23304
rect 17552 23264 17558 23276
rect 19337 23273 19349 23276
rect 19383 23273 19395 23307
rect 19337 23267 19395 23273
rect 26786 23264 26792 23316
rect 26844 23304 26850 23316
rect 27065 23307 27123 23313
rect 27065 23304 27077 23307
rect 26844 23276 27077 23304
rect 26844 23264 26850 23276
rect 27065 23273 27077 23276
rect 27111 23273 27123 23307
rect 27065 23267 27123 23273
rect 27249 23307 27307 23313
rect 27249 23273 27261 23307
rect 27295 23304 27307 23307
rect 27338 23304 27344 23316
rect 27295 23276 27344 23304
rect 27295 23273 27307 23276
rect 27249 23267 27307 23273
rect 27338 23264 27344 23276
rect 27396 23264 27402 23316
rect 29546 23264 29552 23316
rect 29604 23304 29610 23316
rect 29641 23307 29699 23313
rect 29641 23304 29653 23307
rect 29604 23276 29653 23304
rect 29604 23264 29610 23276
rect 29641 23273 29653 23276
rect 29687 23273 29699 23307
rect 29641 23267 29699 23273
rect 15470 23196 15476 23248
rect 15528 23236 15534 23248
rect 15841 23239 15899 23245
rect 15841 23236 15853 23239
rect 15528 23208 15853 23236
rect 15528 23196 15534 23208
rect 15841 23205 15853 23208
rect 15887 23205 15899 23239
rect 30098 23236 30104 23248
rect 15841 23199 15899 23205
rect 30024 23208 30104 23236
rect 15856 23168 15884 23199
rect 15856 23140 16528 23168
rect 16500 23112 16528 23140
rect 1762 23100 1768 23112
rect 1723 23072 1768 23100
rect 1762 23060 1768 23072
rect 1820 23060 1826 23112
rect 2409 23103 2467 23109
rect 2409 23069 2421 23103
rect 2455 23100 2467 23103
rect 2455 23072 6914 23100
rect 2455 23069 2467 23072
rect 2409 23063 2467 23069
rect 6886 23032 6914 23072
rect 14182 23060 14188 23112
rect 14240 23100 14246 23112
rect 14461 23103 14519 23109
rect 14461 23100 14473 23103
rect 14240 23072 14473 23100
rect 14240 23060 14246 23072
rect 14461 23069 14473 23072
rect 14507 23069 14519 23103
rect 14461 23063 14519 23069
rect 14728 23103 14786 23109
rect 14728 23069 14740 23103
rect 14774 23100 14786 23103
rect 15562 23100 15568 23112
rect 14774 23072 15568 23100
rect 14774 23069 14786 23072
rect 14728 23063 14786 23069
rect 15562 23060 15568 23072
rect 15620 23060 15626 23112
rect 16298 23100 16304 23112
rect 16259 23072 16304 23100
rect 16298 23060 16304 23072
rect 16356 23060 16362 23112
rect 16482 23060 16488 23112
rect 16540 23100 16546 23112
rect 19426 23100 19432 23112
rect 16540 23072 16633 23100
rect 19387 23072 19432 23100
rect 16540 23060 16546 23072
rect 19426 23060 19432 23072
rect 19484 23060 19490 23112
rect 21637 23103 21695 23109
rect 21637 23069 21649 23103
rect 21683 23100 21695 23103
rect 22002 23100 22008 23112
rect 21683 23072 22008 23100
rect 21683 23069 21695 23072
rect 21637 23063 21695 23069
rect 22002 23060 22008 23072
rect 22060 23060 22066 23112
rect 22094 23060 22100 23112
rect 22152 23100 22158 23112
rect 24397 23103 24455 23109
rect 22152 23072 22197 23100
rect 22152 23060 22158 23072
rect 24397 23069 24409 23103
rect 24443 23100 24455 23103
rect 25038 23100 25044 23112
rect 24443 23072 25044 23100
rect 24443 23069 24455 23072
rect 24397 23063 24455 23069
rect 25038 23060 25044 23072
rect 25096 23060 25102 23112
rect 28258 23060 28264 23112
rect 28316 23100 28322 23112
rect 28629 23103 28687 23109
rect 28629 23100 28641 23103
rect 28316 23072 28641 23100
rect 28316 23060 28322 23072
rect 28629 23069 28641 23072
rect 28675 23069 28687 23103
rect 28810 23100 28816 23112
rect 28771 23072 28816 23100
rect 28629 23063 28687 23069
rect 28810 23060 28816 23072
rect 28868 23060 28874 23112
rect 28994 23100 29000 23112
rect 28955 23072 29000 23100
rect 28994 23060 29000 23072
rect 29052 23060 29058 23112
rect 29822 23060 29828 23112
rect 29880 23109 29886 23112
rect 30024 23109 30052 23208
rect 30098 23196 30104 23208
rect 30156 23196 30162 23248
rect 33778 23236 33784 23248
rect 33739 23208 33784 23236
rect 33778 23196 33784 23208
rect 33836 23196 33842 23248
rect 37826 23196 37832 23248
rect 37884 23236 37890 23248
rect 37884 23208 38148 23236
rect 37884 23196 37890 23208
rect 37182 23168 37188 23180
rect 37143 23140 37188 23168
rect 37182 23128 37188 23140
rect 37240 23128 37246 23180
rect 37918 23168 37924 23180
rect 37879 23140 37924 23168
rect 37918 23128 37924 23140
rect 37976 23128 37982 23180
rect 38120 23177 38148 23208
rect 38105 23171 38163 23177
rect 38105 23137 38117 23171
rect 38151 23137 38163 23171
rect 38105 23131 38163 23137
rect 29880 23103 29929 23109
rect 29880 23069 29883 23103
rect 29917 23069 29929 23103
rect 29880 23063 29929 23069
rect 30009 23103 30067 23109
rect 30009 23069 30021 23103
rect 30055 23069 30067 23103
rect 30009 23063 30067 23069
rect 29880 23060 29886 23063
rect 30098 23060 30104 23112
rect 30156 23100 30162 23112
rect 30285 23103 30343 23109
rect 30156 23072 30201 23100
rect 30156 23060 30162 23072
rect 30285 23069 30297 23103
rect 30331 23100 30343 23103
rect 30926 23100 30932 23112
rect 30331 23072 30932 23100
rect 30331 23069 30343 23072
rect 30285 23063 30343 23069
rect 30926 23060 30932 23072
rect 30984 23060 30990 23112
rect 32585 23103 32643 23109
rect 32585 23069 32597 23103
rect 32631 23100 32643 23103
rect 32674 23100 32680 23112
rect 32631 23072 32680 23100
rect 32631 23069 32643 23072
rect 32585 23063 32643 23069
rect 32674 23060 32680 23072
rect 32732 23060 32738 23112
rect 33594 23100 33600 23112
rect 33555 23072 33600 23100
rect 33594 23060 33600 23072
rect 33652 23060 33658 23112
rect 35434 23100 35440 23112
rect 35395 23072 35440 23100
rect 35434 23060 35440 23072
rect 35492 23060 35498 23112
rect 9582 23032 9588 23044
rect 6886 23004 9588 23032
rect 9582 22992 9588 23004
rect 9640 23032 9646 23044
rect 14550 23032 14556 23044
rect 9640 23004 14556 23032
rect 9640 22992 9646 23004
rect 14550 22992 14556 23004
rect 14608 22992 14614 23044
rect 24670 23041 24676 23044
rect 24664 22995 24676 23041
rect 24728 23032 24734 23044
rect 27430 23032 27436 23044
rect 24728 23004 24764 23032
rect 27391 23004 27436 23032
rect 24670 22992 24676 22995
rect 24728 22992 24734 23004
rect 27430 22992 27436 23004
rect 27488 22992 27494 23044
rect 28721 23035 28779 23041
rect 28721 23001 28733 23035
rect 28767 23032 28779 23035
rect 28902 23032 28908 23044
rect 28767 23004 28908 23032
rect 28767 23001 28779 23004
rect 28721 22995 28779 23001
rect 28902 22992 28908 23004
rect 28960 23032 28966 23044
rect 28960 23004 29960 23032
rect 28960 22992 28966 23004
rect 1946 22924 1952 22976
rect 2004 22964 2010 22976
rect 2317 22967 2375 22973
rect 2317 22964 2329 22967
rect 2004 22936 2329 22964
rect 2004 22924 2010 22936
rect 2317 22933 2329 22936
rect 2363 22933 2375 22967
rect 2317 22927 2375 22933
rect 20898 22924 20904 22976
rect 20956 22964 20962 22976
rect 21545 22967 21603 22973
rect 21545 22964 21557 22967
rect 20956 22936 21557 22964
rect 20956 22924 20962 22936
rect 21545 22933 21557 22936
rect 21591 22933 21603 22967
rect 21545 22927 21603 22933
rect 21634 22924 21640 22976
rect 21692 22964 21698 22976
rect 22002 22964 22008 22976
rect 21692 22936 22008 22964
rect 21692 22924 21698 22936
rect 22002 22924 22008 22936
rect 22060 22964 22066 22976
rect 22189 22967 22247 22973
rect 22189 22964 22201 22967
rect 22060 22936 22201 22964
rect 22060 22924 22066 22936
rect 22189 22933 22201 22936
rect 22235 22933 22247 22967
rect 25774 22964 25780 22976
rect 25735 22936 25780 22964
rect 22189 22927 22247 22933
rect 25774 22924 25780 22936
rect 25832 22964 25838 22976
rect 26970 22964 26976 22976
rect 25832 22936 26976 22964
rect 25832 22924 25838 22936
rect 26970 22924 26976 22936
rect 27028 22964 27034 22976
rect 27223 22967 27281 22973
rect 27223 22964 27235 22967
rect 27028 22936 27235 22964
rect 27028 22924 27034 22936
rect 27223 22933 27235 22936
rect 27269 22933 27281 22967
rect 27223 22927 27281 22933
rect 28445 22967 28503 22973
rect 28445 22933 28457 22967
rect 28491 22964 28503 22967
rect 29730 22964 29736 22976
rect 28491 22936 29736 22964
rect 28491 22933 28503 22936
rect 28445 22927 28503 22933
rect 29730 22924 29736 22936
rect 29788 22924 29794 22976
rect 29932 22964 29960 23004
rect 32122 22992 32128 23044
rect 32180 23032 32186 23044
rect 32318 23035 32376 23041
rect 32318 23032 32330 23035
rect 32180 23004 32330 23032
rect 32180 22992 32186 23004
rect 32318 23001 32330 23004
rect 32364 23001 32376 23035
rect 32318 22995 32376 23001
rect 31018 22964 31024 22976
rect 29932 22936 31024 22964
rect 31018 22924 31024 22936
rect 31076 22924 31082 22976
rect 31202 22964 31208 22976
rect 31163 22936 31208 22964
rect 31202 22924 31208 22936
rect 31260 22924 31266 22976
rect 35345 22967 35403 22973
rect 35345 22933 35357 22967
rect 35391 22964 35403 22967
rect 35526 22964 35532 22976
rect 35391 22936 35532 22964
rect 35391 22933 35403 22936
rect 35345 22927 35403 22933
rect 35526 22924 35532 22936
rect 35584 22924 35590 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 19245 22763 19303 22769
rect 19245 22729 19257 22763
rect 19291 22760 19303 22763
rect 19426 22760 19432 22772
rect 19291 22732 19432 22760
rect 19291 22729 19303 22732
rect 19245 22723 19303 22729
rect 19426 22720 19432 22732
rect 19484 22720 19490 22772
rect 20806 22720 20812 22772
rect 20864 22760 20870 22772
rect 20993 22763 21051 22769
rect 20993 22760 21005 22763
rect 20864 22732 21005 22760
rect 20864 22720 20870 22732
rect 20993 22729 21005 22732
rect 21039 22729 21051 22763
rect 24670 22760 24676 22772
rect 24631 22732 24676 22760
rect 20993 22723 21051 22729
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 32122 22760 32128 22772
rect 32083 22732 32128 22760
rect 32122 22720 32128 22732
rect 32180 22720 32186 22772
rect 33594 22720 33600 22772
rect 33652 22760 33658 22772
rect 33873 22763 33931 22769
rect 33873 22760 33885 22763
rect 33652 22732 33885 22760
rect 33652 22720 33658 22732
rect 33873 22729 33885 22732
rect 33919 22729 33931 22763
rect 33873 22723 33931 22729
rect 33980 22732 35296 22760
rect 1946 22692 1952 22704
rect 1907 22664 1952 22692
rect 1946 22652 1952 22664
rect 2004 22652 2010 22704
rect 18132 22695 18190 22701
rect 18132 22661 18144 22695
rect 18178 22692 18190 22695
rect 18690 22692 18696 22704
rect 18178 22664 18696 22692
rect 18178 22661 18190 22664
rect 18132 22655 18190 22661
rect 18690 22652 18696 22664
rect 18748 22652 18754 22704
rect 22370 22692 22376 22704
rect 22331 22664 22376 22692
rect 22370 22652 22376 22664
rect 22428 22652 22434 22704
rect 24946 22692 24952 22704
rect 23584 22664 24952 22692
rect 1762 22624 1768 22636
rect 1723 22596 1768 22624
rect 1762 22584 1768 22596
rect 1820 22584 1826 22636
rect 16482 22584 16488 22636
rect 16540 22624 16546 22636
rect 16669 22627 16727 22633
rect 16669 22624 16681 22627
rect 16540 22596 16681 22624
rect 16540 22584 16546 22596
rect 16669 22593 16681 22596
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 20625 22627 20683 22633
rect 20625 22593 20637 22627
rect 20671 22624 20683 22627
rect 21634 22624 21640 22636
rect 20671 22596 21640 22624
rect 20671 22593 20683 22596
rect 20625 22587 20683 22593
rect 21634 22584 21640 22596
rect 21692 22584 21698 22636
rect 23106 22624 23112 22636
rect 23067 22596 23112 22624
rect 23106 22584 23112 22596
rect 23164 22584 23170 22636
rect 23584 22633 23612 22664
rect 24596 22633 24624 22664
rect 24946 22652 24952 22664
rect 25004 22692 25010 22704
rect 25682 22692 25688 22704
rect 25004 22664 25688 22692
rect 25004 22652 25010 22664
rect 25682 22652 25688 22664
rect 25740 22652 25746 22704
rect 28813 22695 28871 22701
rect 28813 22661 28825 22695
rect 28859 22692 28871 22695
rect 28902 22692 28908 22704
rect 28859 22664 28908 22692
rect 28859 22661 28871 22664
rect 28813 22655 28871 22661
rect 28902 22652 28908 22664
rect 28960 22652 28966 22704
rect 32858 22692 32864 22704
rect 32508 22664 32864 22692
rect 23569 22627 23627 22633
rect 23569 22593 23581 22627
rect 23615 22593 23627 22627
rect 23569 22587 23627 22593
rect 23753 22627 23811 22633
rect 23753 22593 23765 22627
rect 23799 22593 23811 22627
rect 23753 22587 23811 22593
rect 24581 22627 24639 22633
rect 24581 22593 24593 22627
rect 24627 22593 24639 22627
rect 24581 22587 24639 22593
rect 24765 22627 24823 22633
rect 24765 22593 24777 22627
rect 24811 22624 24823 22627
rect 25774 22624 25780 22636
rect 24811 22596 25780 22624
rect 24811 22593 24823 22596
rect 24765 22587 24823 22593
rect 2774 22556 2780 22568
rect 2735 22528 2780 22556
rect 2774 22516 2780 22528
rect 2832 22516 2838 22568
rect 17862 22556 17868 22568
rect 17823 22528 17868 22556
rect 17862 22516 17868 22528
rect 17920 22516 17926 22568
rect 20530 22556 20536 22568
rect 20491 22528 20536 22556
rect 20530 22516 20536 22528
rect 20588 22516 20594 22568
rect 23290 22516 23296 22568
rect 23348 22556 23354 22568
rect 23768 22556 23796 22587
rect 25774 22584 25780 22596
rect 25832 22584 25838 22636
rect 28258 22584 28264 22636
rect 28316 22624 28322 22636
rect 28629 22627 28687 22633
rect 28629 22624 28641 22627
rect 28316 22596 28641 22624
rect 28316 22584 28322 22596
rect 28629 22593 28641 22596
rect 28675 22593 28687 22627
rect 28629 22587 28687 22593
rect 28997 22627 29055 22633
rect 28997 22593 29009 22627
rect 29043 22624 29055 22627
rect 29457 22627 29515 22633
rect 29457 22624 29469 22627
rect 29043 22596 29469 22624
rect 29043 22593 29055 22596
rect 28997 22587 29055 22593
rect 29457 22593 29469 22596
rect 29503 22593 29515 22627
rect 29638 22624 29644 22636
rect 29599 22596 29644 22624
rect 29457 22587 29515 22593
rect 29638 22584 29644 22596
rect 29696 22584 29702 22636
rect 29730 22584 29736 22636
rect 29788 22624 29794 22636
rect 30009 22627 30067 22633
rect 29788 22596 29833 22624
rect 29788 22584 29794 22596
rect 30009 22593 30021 22627
rect 30055 22593 30067 22627
rect 30009 22587 30067 22593
rect 23348 22528 23796 22556
rect 23348 22516 23354 22528
rect 29822 22516 29828 22568
rect 29880 22556 29886 22568
rect 29880 22528 29925 22556
rect 29880 22516 29886 22528
rect 29546 22448 29552 22500
rect 29604 22488 29610 22500
rect 30024 22488 30052 22587
rect 30374 22584 30380 22636
rect 30432 22624 30438 22636
rect 31202 22624 31208 22636
rect 30432 22596 31208 22624
rect 30432 22584 30438 22596
rect 31202 22584 31208 22596
rect 31260 22624 31266 22636
rect 32508 22633 32536 22664
rect 32858 22652 32864 22664
rect 32916 22692 32922 22704
rect 33980 22692 34008 22732
rect 32916 22664 34008 22692
rect 34517 22695 34575 22701
rect 32916 22652 32922 22664
rect 34517 22661 34529 22695
rect 34563 22692 34575 22695
rect 34563 22664 35204 22692
rect 34563 22661 34575 22664
rect 34517 22655 34575 22661
rect 32401 22627 32459 22633
rect 32401 22624 32413 22627
rect 31260 22596 32413 22624
rect 31260 22584 31266 22596
rect 32401 22593 32413 22596
rect 32447 22593 32459 22627
rect 32401 22587 32459 22593
rect 32493 22627 32551 22633
rect 32493 22593 32505 22627
rect 32539 22593 32551 22627
rect 32493 22587 32551 22593
rect 32582 22584 32588 22636
rect 32640 22624 32646 22636
rect 32640 22596 32685 22624
rect 32640 22584 32646 22596
rect 32766 22584 32772 22636
rect 32824 22624 32830 22636
rect 35176 22633 35204 22664
rect 35268 22633 35296 22732
rect 34977 22627 35035 22633
rect 34977 22624 34989 22627
rect 32824 22596 34989 22624
rect 32824 22584 32830 22596
rect 34977 22593 34989 22596
rect 35023 22593 35035 22627
rect 34977 22587 35035 22593
rect 35161 22627 35219 22633
rect 35161 22593 35173 22627
rect 35207 22593 35219 22627
rect 35161 22587 35219 22593
rect 35253 22627 35311 22633
rect 35253 22593 35265 22627
rect 35299 22593 35311 22627
rect 35253 22587 35311 22593
rect 35345 22627 35403 22633
rect 35345 22593 35357 22627
rect 35391 22593 35403 22627
rect 36262 22624 36268 22636
rect 36223 22596 36268 22624
rect 35345 22587 35403 22593
rect 34238 22556 34244 22568
rect 34199 22528 34244 22556
rect 34238 22516 34244 22528
rect 34296 22516 34302 22568
rect 34333 22559 34391 22565
rect 34333 22525 34345 22559
rect 34379 22556 34391 22559
rect 34514 22556 34520 22568
rect 34379 22528 34520 22556
rect 34379 22525 34391 22528
rect 34333 22519 34391 22525
rect 34514 22516 34520 22528
rect 34572 22516 34578 22568
rect 35360 22556 35388 22587
rect 36262 22584 36268 22596
rect 36320 22584 36326 22636
rect 36081 22559 36139 22565
rect 36081 22556 36093 22559
rect 34624 22528 36093 22556
rect 34624 22500 34652 22528
rect 36081 22525 36093 22528
rect 36127 22525 36139 22559
rect 36081 22519 36139 22525
rect 34606 22488 34612 22500
rect 29604 22460 34612 22488
rect 29604 22448 29610 22460
rect 34606 22448 34612 22460
rect 34664 22448 34670 22500
rect 16761 22423 16819 22429
rect 16761 22389 16773 22423
rect 16807 22420 16819 22423
rect 16942 22420 16948 22432
rect 16807 22392 16948 22420
rect 16807 22389 16819 22392
rect 16761 22383 16819 22389
rect 16942 22380 16948 22392
rect 17000 22380 17006 22432
rect 22278 22420 22284 22432
rect 22239 22392 22284 22420
rect 22278 22380 22284 22392
rect 22336 22380 22342 22432
rect 22462 22380 22468 22432
rect 22520 22420 22526 22432
rect 23017 22423 23075 22429
rect 23017 22420 23029 22423
rect 22520 22392 23029 22420
rect 22520 22380 22526 22392
rect 23017 22389 23029 22392
rect 23063 22389 23075 22423
rect 23017 22383 23075 22389
rect 23569 22423 23627 22429
rect 23569 22389 23581 22423
rect 23615 22420 23627 22423
rect 24210 22420 24216 22432
rect 23615 22392 24216 22420
rect 23615 22389 23627 22392
rect 23569 22383 23627 22389
rect 24210 22380 24216 22392
rect 24268 22380 24274 22432
rect 30190 22420 30196 22432
rect 30151 22392 30196 22420
rect 30190 22380 30196 22392
rect 30248 22380 30254 22432
rect 35618 22420 35624 22432
rect 35579 22392 35624 22420
rect 35618 22380 35624 22392
rect 35676 22380 35682 22432
rect 37826 22420 37832 22432
rect 37787 22392 37832 22420
rect 37826 22380 37832 22392
rect 37884 22380 37890 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 26605 22219 26663 22225
rect 26605 22185 26617 22219
rect 26651 22216 26663 22219
rect 26786 22216 26792 22228
rect 26651 22188 26792 22216
rect 26651 22185 26663 22188
rect 26605 22179 26663 22185
rect 26786 22176 26792 22188
rect 26844 22176 26850 22228
rect 28258 22216 28264 22228
rect 28219 22188 28264 22216
rect 28258 22176 28264 22188
rect 28316 22176 28322 22228
rect 32217 22219 32275 22225
rect 32217 22185 32229 22219
rect 32263 22216 32275 22219
rect 32582 22216 32588 22228
rect 32263 22188 32588 22216
rect 32263 22185 32275 22188
rect 32217 22179 32275 22185
rect 32582 22176 32588 22188
rect 32640 22176 32646 22228
rect 34149 22219 34207 22225
rect 34149 22185 34161 22219
rect 34195 22216 34207 22219
rect 34238 22216 34244 22228
rect 34195 22188 34244 22216
rect 34195 22185 34207 22188
rect 34149 22179 34207 22185
rect 34238 22176 34244 22188
rect 34296 22176 34302 22228
rect 20714 22148 20720 22160
rect 20675 22120 20720 22148
rect 20714 22108 20720 22120
rect 20772 22108 20778 22160
rect 1854 22080 1860 22092
rect 1815 22052 1860 22080
rect 1854 22040 1860 22052
rect 1912 22040 1918 22092
rect 15746 22080 15752 22092
rect 15707 22052 15752 22080
rect 15746 22040 15752 22052
rect 15804 22040 15810 22092
rect 16114 22040 16120 22092
rect 16172 22080 16178 22092
rect 16393 22083 16451 22089
rect 16393 22080 16405 22083
rect 16172 22052 16405 22080
rect 16172 22040 16178 22052
rect 16393 22049 16405 22052
rect 16439 22049 16451 22083
rect 16393 22043 16451 22049
rect 16482 22040 16488 22092
rect 16540 22080 16546 22092
rect 16853 22083 16911 22089
rect 16853 22080 16865 22083
rect 16540 22052 16865 22080
rect 16540 22040 16546 22052
rect 16853 22049 16865 22052
rect 16899 22049 16911 22083
rect 16853 22043 16911 22049
rect 20441 22083 20499 22089
rect 20441 22049 20453 22083
rect 20487 22080 20499 22083
rect 20530 22080 20536 22092
rect 20487 22052 20536 22080
rect 20487 22049 20499 22052
rect 20441 22043 20499 22049
rect 20530 22040 20536 22052
rect 20588 22040 20594 22092
rect 26694 22040 26700 22092
rect 26752 22080 26758 22092
rect 26789 22083 26847 22089
rect 26789 22080 26801 22083
rect 26752 22052 26801 22080
rect 26752 22040 26758 22052
rect 26789 22049 26801 22052
rect 26835 22049 26847 22083
rect 34422 22080 34428 22092
rect 26789 22043 26847 22049
rect 33796 22052 34428 22080
rect 1394 22012 1400 22024
rect 1355 21984 1400 22012
rect 1394 21972 1400 21984
rect 1452 21972 1458 22024
rect 15654 22012 15660 22024
rect 15615 21984 15660 22012
rect 15654 21972 15660 21984
rect 15712 22012 15718 22024
rect 15838 22012 15844 22024
rect 15712 21984 15844 22012
rect 15712 21972 15718 21984
rect 15838 21972 15844 21984
rect 15896 21972 15902 22024
rect 16574 22012 16580 22024
rect 16535 21984 16580 22012
rect 16574 21972 16580 21984
rect 16632 21972 16638 22024
rect 16666 21972 16672 22024
rect 16724 22012 16730 22024
rect 16942 22012 16948 22024
rect 16724 21984 16948 22012
rect 16724 21972 16730 21984
rect 16942 21972 16948 21984
rect 17000 21972 17006 22024
rect 20349 22015 20407 22021
rect 20349 21981 20361 22015
rect 20395 22012 20407 22015
rect 20714 22012 20720 22024
rect 20395 21984 20720 22012
rect 20395 21981 20407 21984
rect 20349 21975 20407 21981
rect 20714 21972 20720 21984
rect 20772 21972 20778 22024
rect 22370 22012 22376 22024
rect 22331 21984 22376 22012
rect 22370 21972 22376 21984
rect 22428 21972 22434 22024
rect 22462 21972 22468 22024
rect 22520 22012 22526 22024
rect 22646 22012 22652 22024
rect 22520 21984 22565 22012
rect 22607 21984 22652 22012
rect 22520 21972 22526 21984
rect 22646 21972 22652 21984
rect 22704 21972 22710 22024
rect 22741 22015 22799 22021
rect 22741 21981 22753 22015
rect 22787 22012 22799 22015
rect 23293 22015 23351 22021
rect 23293 22012 23305 22015
rect 22787 21984 23305 22012
rect 22787 21981 22799 21984
rect 22741 21975 22799 21981
rect 23293 21981 23305 21984
rect 23339 21981 23351 22015
rect 23293 21975 23351 21981
rect 23382 21972 23388 22024
rect 23440 22012 23446 22024
rect 26513 22015 26571 22021
rect 23440 21984 23485 22012
rect 23440 21972 23446 21984
rect 26513 21981 26525 22015
rect 26559 21981 26571 22015
rect 26513 21975 26571 21981
rect 28169 22015 28227 22021
rect 28169 21981 28181 22015
rect 28215 21981 28227 22015
rect 32122 22012 32128 22024
rect 32083 21984 32128 22012
rect 28169 21975 28227 21981
rect 1581 21947 1639 21953
rect 1581 21913 1593 21947
rect 1627 21944 1639 21947
rect 2038 21944 2044 21956
rect 1627 21916 2044 21944
rect 1627 21913 1639 21916
rect 1581 21907 1639 21913
rect 2038 21904 2044 21916
rect 2096 21904 2102 21956
rect 26418 21904 26424 21956
rect 26476 21944 26482 21956
rect 26528 21944 26556 21975
rect 28184 21944 28212 21975
rect 32122 21972 32128 21984
rect 32180 21972 32186 22024
rect 32214 21972 32220 22024
rect 32272 22012 32278 22024
rect 32309 22015 32367 22021
rect 32309 22012 32321 22015
rect 32272 21984 32321 22012
rect 32272 21972 32278 21984
rect 32309 21981 32321 21984
rect 32355 22012 32367 22015
rect 33686 22012 33692 22024
rect 32355 21984 33692 22012
rect 32355 21981 32367 21984
rect 32309 21975 32367 21981
rect 33686 21972 33692 21984
rect 33744 21972 33750 22024
rect 33796 22021 33824 22052
rect 34422 22040 34428 22052
rect 34480 22080 34486 22092
rect 35253 22083 35311 22089
rect 35253 22080 35265 22083
rect 34480 22052 35265 22080
rect 34480 22040 34486 22052
rect 35253 22049 35265 22052
rect 35299 22049 35311 22083
rect 35526 22080 35532 22092
rect 35487 22052 35532 22080
rect 35253 22043 35311 22049
rect 35526 22040 35532 22052
rect 35584 22040 35590 22092
rect 37182 22080 37188 22092
rect 37143 22052 37188 22080
rect 37182 22040 37188 22052
rect 37240 22040 37246 22092
rect 37826 22040 37832 22092
rect 37884 22080 37890 22092
rect 38105 22083 38163 22089
rect 38105 22080 38117 22083
rect 37884 22052 38117 22080
rect 37884 22040 37890 22052
rect 38105 22049 38117 22052
rect 38151 22049 38163 22083
rect 38105 22043 38163 22049
rect 33781 22015 33839 22021
rect 33781 21981 33793 22015
rect 33827 21981 33839 22015
rect 33781 21975 33839 21981
rect 33965 22015 34023 22021
rect 33965 21981 33977 22015
rect 34011 22012 34023 22015
rect 34790 22012 34796 22024
rect 34011 21984 34796 22012
rect 34011 21981 34023 21984
rect 33965 21975 34023 21981
rect 34790 21972 34796 21984
rect 34848 21972 34854 22024
rect 35621 22015 35679 22021
rect 35621 21981 35633 22015
rect 35667 22012 35679 22015
rect 36262 22012 36268 22024
rect 35667 21984 36268 22012
rect 35667 21981 35679 21984
rect 35621 21975 35679 21981
rect 36262 21972 36268 21984
rect 36320 21972 36326 22024
rect 26476 21916 28212 21944
rect 26476 21904 26482 21916
rect 37458 21904 37464 21956
rect 37516 21944 37522 21956
rect 37921 21947 37979 21953
rect 37921 21944 37933 21947
rect 37516 21916 37933 21944
rect 37516 21904 37522 21916
rect 37921 21913 37933 21916
rect 37967 21913 37979 21947
rect 37921 21907 37979 21913
rect 22189 21879 22247 21885
rect 22189 21845 22201 21879
rect 22235 21876 22247 21879
rect 22554 21876 22560 21888
rect 22235 21848 22560 21876
rect 22235 21845 22247 21848
rect 22189 21839 22247 21845
rect 22554 21836 22560 21848
rect 22612 21836 22618 21888
rect 26789 21879 26847 21885
rect 26789 21845 26801 21879
rect 26835 21876 26847 21879
rect 27798 21876 27804 21888
rect 26835 21848 27804 21876
rect 26835 21845 26847 21848
rect 26789 21839 26847 21845
rect 27798 21836 27804 21848
rect 27856 21836 27862 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 2038 21672 2044 21684
rect 1999 21644 2044 21672
rect 2038 21632 2044 21644
rect 2096 21632 2102 21684
rect 16574 21632 16580 21684
rect 16632 21672 16638 21684
rect 17037 21675 17095 21681
rect 17037 21672 17049 21675
rect 16632 21644 17049 21672
rect 16632 21632 16638 21644
rect 17037 21641 17049 21644
rect 17083 21641 17095 21675
rect 18046 21672 18052 21684
rect 17037 21635 17095 21641
rect 17420 21644 18052 21672
rect 15194 21604 15200 21616
rect 6886 21576 15200 21604
rect 2133 21539 2191 21545
rect 2133 21505 2145 21539
rect 2179 21536 2191 21539
rect 2406 21536 2412 21548
rect 2179 21508 2412 21536
rect 2179 21505 2191 21508
rect 2133 21499 2191 21505
rect 2406 21496 2412 21508
rect 2464 21536 2470 21548
rect 6886 21536 6914 21576
rect 15194 21564 15200 21576
rect 15252 21564 15258 21616
rect 16206 21564 16212 21616
rect 16264 21604 16270 21616
rect 17420 21613 17448 21644
rect 18046 21632 18052 21644
rect 18104 21672 18110 21684
rect 19521 21675 19579 21681
rect 18104 21644 18736 21672
rect 18104 21632 18110 21644
rect 17313 21607 17371 21613
rect 17313 21604 17325 21607
rect 16264 21576 17325 21604
rect 16264 21564 16270 21576
rect 17313 21573 17325 21576
rect 17359 21573 17371 21607
rect 17313 21567 17371 21573
rect 17405 21607 17463 21613
rect 17405 21573 17417 21607
rect 17451 21573 17463 21607
rect 17405 21567 17463 21573
rect 2464 21508 6914 21536
rect 2464 21496 2470 21508
rect 7834 21496 7840 21548
rect 7892 21536 7898 21548
rect 7929 21539 7987 21545
rect 7929 21536 7941 21539
rect 7892 21508 7941 21536
rect 7892 21496 7898 21508
rect 7929 21505 7941 21508
rect 7975 21505 7987 21539
rect 7929 21499 7987 21505
rect 17216 21539 17274 21545
rect 17216 21505 17228 21539
rect 17262 21536 17274 21539
rect 17262 21508 17356 21536
rect 17262 21505 17274 21508
rect 17216 21499 17274 21505
rect 8754 21468 8760 21480
rect 8715 21440 8760 21468
rect 8754 21428 8760 21440
rect 8812 21428 8818 21480
rect 17328 21468 17356 21508
rect 17494 21496 17500 21548
rect 17552 21536 17558 21548
rect 18708 21545 18736 21644
rect 19521 21641 19533 21675
rect 19567 21641 19579 21675
rect 19521 21635 19579 21641
rect 20625 21675 20683 21681
rect 20625 21641 20637 21675
rect 20671 21641 20683 21675
rect 20625 21635 20683 21641
rect 19334 21604 19340 21616
rect 18892 21576 19340 21604
rect 18892 21545 18920 21576
rect 19334 21564 19340 21576
rect 19392 21564 19398 21616
rect 17588 21539 17646 21545
rect 17588 21536 17600 21539
rect 17552 21508 17600 21536
rect 17552 21496 17558 21508
rect 17588 21505 17600 21508
rect 17634 21505 17646 21539
rect 17588 21499 17646 21505
rect 17681 21539 17739 21545
rect 17681 21505 17693 21539
rect 17727 21536 17739 21539
rect 18325 21539 18383 21545
rect 18325 21536 18337 21539
rect 17727 21508 18337 21536
rect 17727 21505 17739 21508
rect 17681 21499 17739 21505
rect 18325 21505 18337 21508
rect 18371 21505 18383 21539
rect 18325 21499 18383 21505
rect 18509 21539 18567 21545
rect 18509 21505 18521 21539
rect 18555 21505 18567 21539
rect 18509 21499 18567 21505
rect 18693 21539 18751 21545
rect 18693 21505 18705 21539
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 18877 21539 18935 21545
rect 18877 21505 18889 21539
rect 18923 21505 18935 21539
rect 18877 21499 18935 21505
rect 19061 21539 19119 21545
rect 19061 21505 19073 21539
rect 19107 21536 19119 21539
rect 19536 21536 19564 21635
rect 19107 21508 19564 21536
rect 19107 21505 19119 21508
rect 19061 21499 19119 21505
rect 17604 21468 17632 21499
rect 18524 21468 18552 21499
rect 19610 21496 19616 21548
rect 19668 21536 19674 21548
rect 19705 21539 19763 21545
rect 19705 21536 19717 21539
rect 19668 21508 19717 21536
rect 19668 21496 19674 21508
rect 19705 21505 19717 21508
rect 19751 21505 19763 21539
rect 19705 21499 19763 21505
rect 19797 21539 19855 21545
rect 19797 21505 19809 21539
rect 19843 21505 19855 21539
rect 19797 21499 19855 21505
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21536 19947 21539
rect 19978 21536 19984 21548
rect 19935 21508 19984 21536
rect 19935 21505 19947 21508
rect 19889 21499 19947 21505
rect 17328 21440 17540 21468
rect 17604 21440 18552 21468
rect 18785 21471 18843 21477
rect 17512 21412 17540 21440
rect 18785 21437 18797 21471
rect 18831 21468 18843 21471
rect 19150 21468 19156 21480
rect 18831 21440 19156 21468
rect 18831 21437 18843 21440
rect 18785 21431 18843 21437
rect 19150 21428 19156 21440
rect 19208 21468 19214 21480
rect 19812 21468 19840 21499
rect 19978 21496 19984 21508
rect 20036 21496 20042 21548
rect 20073 21539 20131 21545
rect 20073 21505 20085 21539
rect 20119 21536 20131 21539
rect 20640 21536 20668 21635
rect 20714 21632 20720 21684
rect 20772 21672 20778 21684
rect 20772 21644 20944 21672
rect 20772 21632 20778 21644
rect 20916 21613 20944 21644
rect 22646 21632 22652 21684
rect 22704 21672 22710 21684
rect 23109 21675 23167 21681
rect 23109 21672 23121 21675
rect 22704 21644 23121 21672
rect 22704 21632 22710 21644
rect 23109 21641 23121 21644
rect 23155 21641 23167 21675
rect 26418 21672 26424 21684
rect 26379 21644 26424 21672
rect 23109 21635 23167 21641
rect 26418 21632 26424 21644
rect 26476 21632 26482 21684
rect 30466 21672 30472 21684
rect 28460 21644 30472 21672
rect 20901 21607 20959 21613
rect 20901 21573 20913 21607
rect 20947 21573 20959 21607
rect 20901 21567 20959 21573
rect 21192 21576 22048 21604
rect 21192 21545 21220 21576
rect 22020 21548 22048 21576
rect 22278 21564 22284 21616
rect 22336 21604 22342 21616
rect 25308 21607 25366 21613
rect 22336 21576 24532 21604
rect 22336 21564 22342 21576
rect 20119 21508 20668 21536
rect 20804 21539 20862 21545
rect 20119 21505 20131 21508
rect 20073 21499 20131 21505
rect 20804 21505 20816 21539
rect 20850 21505 20862 21539
rect 20804 21499 20862 21505
rect 20993 21539 21051 21545
rect 20993 21505 21005 21539
rect 21039 21505 21051 21539
rect 20993 21499 21051 21505
rect 21176 21539 21234 21545
rect 21176 21505 21188 21539
rect 21222 21505 21234 21539
rect 21176 21499 21234 21505
rect 21269 21539 21327 21545
rect 21269 21505 21281 21539
rect 21315 21536 21327 21539
rect 21821 21539 21879 21545
rect 21821 21536 21833 21539
rect 21315 21508 21833 21536
rect 21315 21505 21327 21508
rect 21269 21499 21327 21505
rect 21821 21505 21833 21508
rect 21867 21505 21879 21539
rect 22002 21536 22008 21548
rect 21963 21508 22008 21536
rect 21821 21499 21879 21505
rect 19208 21440 19840 21468
rect 19208 21428 19214 21440
rect 20346 21428 20352 21480
rect 20404 21468 20410 21480
rect 20824 21468 20852 21499
rect 20404 21440 20852 21468
rect 21008 21468 21036 21499
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 22094 21496 22100 21548
rect 22152 21536 22158 21548
rect 22373 21539 22431 21545
rect 22373 21536 22385 21539
rect 22152 21508 22385 21536
rect 22152 21496 22158 21508
rect 22373 21505 22385 21508
rect 22419 21505 22431 21539
rect 22554 21536 22560 21548
rect 22515 21508 22560 21536
rect 22373 21499 22431 21505
rect 22554 21496 22560 21508
rect 22612 21496 22618 21548
rect 24210 21496 24216 21548
rect 24268 21545 24274 21548
rect 24504 21545 24532 21576
rect 25308 21573 25320 21607
rect 25354 21604 25366 21607
rect 27893 21607 27951 21613
rect 27893 21604 27905 21607
rect 25354 21576 27905 21604
rect 25354 21573 25366 21576
rect 25308 21567 25366 21573
rect 27893 21573 27905 21576
rect 27939 21573 27951 21607
rect 27893 21567 27951 21573
rect 24268 21536 24280 21545
rect 24489 21539 24547 21545
rect 24268 21508 24313 21536
rect 24268 21499 24280 21508
rect 24489 21505 24501 21539
rect 24535 21536 24547 21539
rect 25038 21536 25044 21548
rect 24535 21508 25044 21536
rect 24535 21505 24547 21508
rect 24489 21499 24547 21505
rect 24268 21496 24274 21499
rect 25038 21496 25044 21508
rect 25096 21496 25102 21548
rect 26418 21496 26424 21548
rect 26476 21536 26482 21548
rect 26970 21536 26976 21548
rect 26476 21508 26976 21536
rect 26476 21496 26482 21508
rect 26970 21496 26976 21508
rect 27028 21496 27034 21548
rect 27157 21539 27215 21545
rect 27157 21505 27169 21539
rect 27203 21505 27215 21539
rect 27798 21536 27804 21548
rect 27759 21508 27804 21536
rect 27157 21499 27215 21505
rect 22189 21471 22247 21477
rect 22189 21468 22201 21471
rect 21008 21440 22201 21468
rect 20404 21428 20410 21440
rect 22189 21437 22201 21440
rect 22235 21437 22247 21471
rect 22189 21431 22247 21437
rect 22281 21471 22339 21477
rect 22281 21437 22293 21471
rect 22327 21468 22339 21471
rect 22462 21468 22468 21480
rect 22327 21440 22468 21468
rect 22327 21437 22339 21440
rect 22281 21431 22339 21437
rect 17494 21360 17500 21412
rect 17552 21360 17558 21412
rect 22204 21400 22232 21431
rect 22462 21428 22468 21440
rect 22520 21428 22526 21480
rect 26786 21428 26792 21480
rect 26844 21468 26850 21480
rect 27172 21468 27200 21499
rect 27798 21496 27804 21508
rect 27856 21496 27862 21548
rect 28460 21545 28488 21644
rect 30466 21632 30472 21644
rect 30524 21672 30530 21684
rect 32122 21672 32128 21684
rect 30524 21644 30788 21672
rect 32083 21644 32128 21672
rect 30524 21632 30530 21644
rect 29733 21607 29791 21613
rect 29733 21573 29745 21607
rect 29779 21604 29791 21607
rect 30760 21604 30788 21644
rect 32122 21632 32128 21644
rect 32180 21632 32186 21684
rect 34514 21672 34520 21684
rect 34475 21644 34520 21672
rect 34514 21632 34520 21644
rect 34572 21632 34578 21684
rect 34624 21644 35894 21672
rect 34624 21604 34652 21644
rect 29779 21576 30696 21604
rect 30760 21576 34652 21604
rect 29779 21573 29791 21576
rect 29733 21567 29791 21573
rect 27985 21539 28043 21545
rect 27985 21505 27997 21539
rect 28031 21505 28043 21539
rect 27985 21499 28043 21505
rect 28445 21539 28503 21545
rect 28445 21505 28457 21539
rect 28491 21505 28503 21539
rect 28445 21499 28503 21505
rect 29641 21539 29699 21545
rect 29641 21505 29653 21539
rect 29687 21536 29699 21539
rect 30098 21536 30104 21548
rect 29687 21508 30104 21536
rect 29687 21505 29699 21508
rect 29641 21499 29699 21505
rect 28000 21468 28028 21499
rect 30098 21496 30104 21508
rect 30156 21496 30162 21548
rect 30285 21539 30343 21545
rect 30285 21505 30297 21539
rect 30331 21536 30343 21539
rect 30374 21536 30380 21548
rect 30331 21508 30380 21536
rect 30331 21505 30343 21508
rect 30285 21499 30343 21505
rect 30374 21496 30380 21508
rect 30432 21496 30438 21548
rect 30668 21545 30696 21576
rect 30469 21539 30527 21545
rect 30469 21505 30481 21539
rect 30515 21505 30527 21539
rect 30469 21499 30527 21505
rect 30561 21539 30619 21545
rect 30561 21505 30573 21539
rect 30607 21505 30619 21539
rect 30561 21499 30619 21505
rect 30653 21539 30711 21545
rect 30653 21505 30665 21539
rect 30699 21536 30711 21539
rect 31478 21536 31484 21548
rect 30699 21508 31484 21536
rect 30699 21505 30711 21508
rect 30653 21499 30711 21505
rect 30484 21468 30512 21499
rect 26844 21440 27200 21468
rect 27356 21440 28028 21468
rect 30300 21440 30512 21468
rect 30576 21468 30604 21499
rect 31478 21496 31484 21508
rect 31536 21496 31542 21548
rect 32493 21539 32551 21545
rect 32493 21505 32505 21539
rect 32539 21505 32551 21539
rect 32493 21499 32551 21505
rect 30834 21468 30840 21480
rect 30576 21440 30840 21468
rect 26844 21428 26850 21440
rect 22922 21400 22928 21412
rect 22204 21372 22928 21400
rect 22922 21360 22928 21372
rect 22980 21360 22986 21412
rect 26510 21292 26516 21344
rect 26568 21332 26574 21344
rect 27356 21341 27384 21440
rect 30300 21412 30328 21440
rect 30834 21428 30840 21440
rect 30892 21428 30898 21480
rect 32401 21471 32459 21477
rect 32401 21437 32413 21471
rect 32447 21437 32459 21471
rect 32508 21468 32536 21499
rect 33042 21496 33048 21548
rect 33100 21536 33106 21548
rect 33137 21539 33195 21545
rect 33137 21536 33149 21539
rect 33100 21508 33149 21536
rect 33100 21496 33106 21508
rect 33137 21505 33149 21508
rect 33183 21505 33195 21539
rect 33318 21536 33324 21548
rect 33279 21508 33324 21536
rect 33137 21499 33195 21505
rect 33318 21496 33324 21508
rect 33376 21496 33382 21548
rect 34422 21536 34428 21548
rect 34383 21508 34428 21536
rect 34422 21496 34428 21508
rect 34480 21496 34486 21548
rect 34609 21539 34667 21545
rect 34609 21505 34621 21539
rect 34655 21536 34667 21539
rect 34790 21536 34796 21548
rect 34655 21508 34796 21536
rect 34655 21505 34667 21508
rect 34609 21499 34667 21505
rect 34790 21496 34796 21508
rect 34848 21496 34854 21548
rect 35069 21539 35127 21545
rect 35069 21505 35081 21539
rect 35115 21536 35127 21539
rect 35158 21536 35164 21548
rect 35115 21508 35164 21536
rect 35115 21505 35127 21508
rect 35069 21499 35127 21505
rect 35158 21496 35164 21508
rect 35216 21496 35222 21548
rect 35336 21539 35394 21545
rect 35336 21505 35348 21539
rect 35382 21536 35394 21539
rect 35618 21536 35624 21548
rect 35382 21508 35624 21536
rect 35382 21505 35394 21508
rect 35336 21499 35394 21505
rect 35618 21496 35624 21508
rect 35676 21496 35682 21548
rect 35866 21536 35894 21644
rect 36262 21632 36268 21684
rect 36320 21672 36326 21684
rect 36449 21675 36507 21681
rect 36449 21672 36461 21675
rect 36320 21644 36461 21672
rect 36320 21632 36326 21644
rect 36449 21641 36461 21644
rect 36495 21641 36507 21675
rect 37458 21672 37464 21684
rect 37419 21644 37464 21672
rect 36449 21635 36507 21641
rect 37458 21632 37464 21644
rect 37516 21632 37522 21684
rect 37369 21539 37427 21545
rect 35866 21508 36952 21536
rect 32582 21468 32588 21480
rect 32508 21440 32588 21468
rect 32401 21431 32459 21437
rect 30282 21360 30288 21412
rect 30340 21360 30346 21412
rect 31202 21360 31208 21412
rect 31260 21400 31266 21412
rect 32416 21400 32444 21431
rect 32582 21428 32588 21440
rect 32640 21468 32646 21480
rect 33229 21471 33287 21477
rect 33229 21468 33241 21471
rect 32640 21440 33241 21468
rect 32640 21428 32646 21440
rect 33229 21437 33241 21440
rect 33275 21437 33287 21471
rect 36924 21468 36952 21508
rect 37369 21505 37381 21539
rect 37415 21536 37427 21539
rect 37642 21536 37648 21548
rect 37415 21508 37648 21536
rect 37415 21505 37427 21508
rect 37369 21499 37427 21505
rect 37642 21496 37648 21508
rect 37700 21496 37706 21548
rect 37826 21468 37832 21480
rect 36924 21440 37832 21468
rect 33229 21431 33287 21437
rect 37826 21428 37832 21440
rect 37884 21428 37890 21480
rect 32766 21400 32772 21412
rect 31260 21372 31524 21400
rect 32416 21372 32772 21400
rect 31260 21360 31266 21372
rect 27341 21335 27399 21341
rect 27341 21332 27353 21335
rect 26568 21304 27353 21332
rect 26568 21292 26574 21304
rect 27341 21301 27353 21304
rect 27387 21301 27399 21335
rect 27341 21295 27399 21301
rect 28629 21335 28687 21341
rect 28629 21301 28641 21335
rect 28675 21332 28687 21335
rect 29086 21332 29092 21344
rect 28675 21304 29092 21332
rect 28675 21301 28687 21304
rect 28629 21295 28687 21301
rect 29086 21292 29092 21304
rect 29144 21292 29150 21344
rect 30837 21335 30895 21341
rect 30837 21301 30849 21335
rect 30883 21332 30895 21335
rect 31386 21332 31392 21344
rect 30883 21304 31392 21332
rect 30883 21301 30895 21304
rect 30837 21295 30895 21301
rect 31386 21292 31392 21304
rect 31444 21292 31450 21344
rect 31496 21332 31524 21372
rect 32766 21360 32772 21372
rect 32824 21360 32830 21412
rect 33134 21332 33140 21344
rect 31496 21304 33140 21332
rect 33134 21292 33140 21304
rect 33192 21292 33198 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1394 21088 1400 21140
rect 1452 21128 1458 21140
rect 1673 21131 1731 21137
rect 1673 21128 1685 21131
rect 1452 21100 1685 21128
rect 1452 21088 1458 21100
rect 1673 21097 1685 21100
rect 1719 21097 1731 21131
rect 16114 21128 16120 21140
rect 16075 21100 16120 21128
rect 1673 21091 1731 21097
rect 16114 21088 16120 21100
rect 16172 21088 16178 21140
rect 16482 21088 16488 21140
rect 16540 21128 16546 21140
rect 16577 21131 16635 21137
rect 16577 21128 16589 21131
rect 16540 21100 16589 21128
rect 16540 21088 16546 21100
rect 16577 21097 16589 21100
rect 16623 21097 16635 21131
rect 19978 21128 19984 21140
rect 19939 21100 19984 21128
rect 16577 21091 16635 21097
rect 19978 21088 19984 21100
rect 20036 21088 20042 21140
rect 26510 21128 26516 21140
rect 26471 21100 26516 21128
rect 26510 21088 26516 21100
rect 26568 21088 26574 21140
rect 26970 21088 26976 21140
rect 27028 21128 27034 21140
rect 27341 21131 27399 21137
rect 27341 21128 27353 21131
rect 27028 21100 27353 21128
rect 27028 21088 27034 21100
rect 27341 21097 27353 21100
rect 27387 21097 27399 21131
rect 27341 21091 27399 21097
rect 28445 21131 28503 21137
rect 28445 21097 28457 21131
rect 28491 21128 28503 21131
rect 29822 21128 29828 21140
rect 28491 21100 29828 21128
rect 28491 21097 28503 21100
rect 28445 21091 28503 21097
rect 29822 21088 29828 21100
rect 29880 21088 29886 21140
rect 31849 21131 31907 21137
rect 31849 21097 31861 21131
rect 31895 21128 31907 21131
rect 31938 21128 31944 21140
rect 31895 21100 31944 21128
rect 31895 21097 31907 21100
rect 31849 21091 31907 21097
rect 31938 21088 31944 21100
rect 31996 21088 32002 21140
rect 9861 21063 9919 21069
rect 9861 21029 9873 21063
rect 9907 21060 9919 21063
rect 9907 21032 35894 21060
rect 9907 21029 9919 21032
rect 9861 21023 9919 21029
rect 8202 20992 8208 21004
rect 8163 20964 8208 20992
rect 8202 20952 8208 20964
rect 8260 20952 8266 21004
rect 16206 20952 16212 21004
rect 16264 20992 16270 21004
rect 16264 20964 16436 20992
rect 16264 20952 16270 20964
rect 7834 20884 7840 20936
rect 7892 20924 7898 20936
rect 7929 20927 7987 20933
rect 7929 20924 7941 20927
rect 7892 20896 7941 20924
rect 7892 20884 7898 20896
rect 7929 20893 7941 20896
rect 7975 20893 7987 20927
rect 8220 20924 8248 20952
rect 16408 20933 16436 20964
rect 22646 20952 22652 21004
rect 22704 20992 22710 21004
rect 23017 20995 23075 21001
rect 23017 20992 23029 20995
rect 22704 20964 23029 20992
rect 22704 20952 22710 20964
rect 23017 20961 23029 20964
rect 23063 20961 23075 20995
rect 23290 20992 23296 21004
rect 23251 20964 23296 20992
rect 23017 20955 23075 20961
rect 23290 20952 23296 20964
rect 23348 20952 23354 21004
rect 26694 20992 26700 21004
rect 26655 20964 26700 20992
rect 26694 20952 26700 20964
rect 26752 20952 26758 21004
rect 30006 20952 30012 21004
rect 30064 20992 30070 21004
rect 30193 20995 30251 21001
rect 30193 20992 30205 20995
rect 30064 20964 30205 20992
rect 30064 20952 30070 20964
rect 30193 20961 30205 20964
rect 30239 20961 30251 20995
rect 30193 20955 30251 20961
rect 30374 20952 30380 21004
rect 30432 20992 30438 21004
rect 31386 20992 31392 21004
rect 30432 20964 30512 20992
rect 31347 20964 31392 20992
rect 30432 20952 30438 20964
rect 9769 20927 9827 20933
rect 9769 20924 9781 20927
rect 8220 20896 9781 20924
rect 7929 20887 7987 20893
rect 9769 20893 9781 20896
rect 9815 20893 9827 20927
rect 9769 20887 9827 20893
rect 16301 20927 16359 20933
rect 16301 20893 16313 20927
rect 16347 20893 16359 20927
rect 16301 20887 16359 20893
rect 16393 20927 16451 20933
rect 16393 20893 16405 20927
rect 16439 20893 16451 20927
rect 16666 20924 16672 20936
rect 16627 20896 16672 20924
rect 16393 20887 16451 20893
rect 16316 20856 16344 20887
rect 16666 20884 16672 20896
rect 16724 20884 16730 20936
rect 20165 20927 20223 20933
rect 20165 20893 20177 20927
rect 20211 20924 20223 20927
rect 20714 20924 20720 20936
rect 20211 20896 20720 20924
rect 20211 20893 20223 20896
rect 20165 20887 20223 20893
rect 20714 20884 20720 20896
rect 20772 20884 20778 20936
rect 26418 20924 26424 20936
rect 26331 20896 26424 20924
rect 26418 20884 26424 20896
rect 26476 20924 26482 20936
rect 28353 20927 28411 20933
rect 28353 20924 28365 20927
rect 26476 20896 28365 20924
rect 26476 20884 26482 20896
rect 17494 20856 17500 20868
rect 16316 20828 17500 20856
rect 17494 20816 17500 20828
rect 17552 20816 17558 20868
rect 20346 20856 20352 20868
rect 20307 20828 20352 20856
rect 20346 20816 20352 20828
rect 20404 20816 20410 20868
rect 26786 20816 26792 20868
rect 26844 20856 26850 20868
rect 27540 20865 27568 20896
rect 28353 20893 28365 20896
rect 28399 20893 28411 20927
rect 29914 20924 29920 20936
rect 29875 20896 29920 20924
rect 28353 20887 28411 20893
rect 29914 20884 29920 20896
rect 29972 20884 29978 20936
rect 30101 20927 30159 20933
rect 30101 20893 30113 20927
rect 30147 20893 30159 20927
rect 30101 20887 30159 20893
rect 27309 20859 27367 20865
rect 27309 20856 27321 20859
rect 26844 20828 27321 20856
rect 26844 20816 26850 20828
rect 27309 20825 27321 20828
rect 27355 20825 27367 20859
rect 27309 20819 27367 20825
rect 27525 20859 27583 20865
rect 27525 20825 27537 20859
rect 27571 20825 27583 20859
rect 27525 20819 27583 20825
rect 29730 20816 29736 20868
rect 29788 20856 29794 20868
rect 30116 20856 30144 20887
rect 30282 20884 30288 20936
rect 30340 20924 30346 20936
rect 30484 20933 30512 20964
rect 31386 20952 31392 20964
rect 31444 20952 31450 21004
rect 31478 20952 31484 21004
rect 31536 20992 31542 21004
rect 33597 20995 33655 21001
rect 31536 20964 31581 20992
rect 31536 20952 31542 20964
rect 33597 20961 33609 20995
rect 33643 20961 33655 20995
rect 33597 20955 33655 20961
rect 33873 20995 33931 21001
rect 33873 20961 33885 20995
rect 33919 20992 33931 20995
rect 34422 20992 34428 21004
rect 33919 20964 34428 20992
rect 33919 20961 33931 20964
rect 33873 20955 33931 20961
rect 30469 20927 30527 20933
rect 30340 20896 30385 20924
rect 30340 20884 30346 20896
rect 30469 20893 30481 20927
rect 30515 20893 30527 20927
rect 30469 20887 30527 20893
rect 31113 20927 31171 20933
rect 31113 20893 31125 20927
rect 31159 20924 31171 20927
rect 31202 20924 31208 20936
rect 31159 20896 31208 20924
rect 31159 20893 31171 20896
rect 31113 20887 31171 20893
rect 31202 20884 31208 20896
rect 31260 20884 31266 20936
rect 31297 20927 31355 20933
rect 31297 20893 31309 20927
rect 31343 20893 31355 20927
rect 31665 20927 31723 20933
rect 31665 20924 31677 20927
rect 31297 20887 31355 20893
rect 31404 20896 31677 20924
rect 29788 20828 30144 20856
rect 30653 20859 30711 20865
rect 29788 20816 29794 20828
rect 30653 20825 30665 20859
rect 30699 20856 30711 20859
rect 31312 20856 31340 20887
rect 30699 20828 31340 20856
rect 30699 20825 30711 20828
rect 30653 20819 30711 20825
rect 26697 20791 26755 20797
rect 26697 20757 26709 20791
rect 26743 20788 26755 20791
rect 26970 20788 26976 20800
rect 26743 20760 26976 20788
rect 26743 20757 26755 20760
rect 26697 20751 26755 20757
rect 26970 20748 26976 20760
rect 27028 20748 27034 20800
rect 27154 20788 27160 20800
rect 27115 20760 27160 20788
rect 27154 20748 27160 20760
rect 27212 20748 27218 20800
rect 30834 20748 30840 20800
rect 30892 20788 30898 20800
rect 31404 20788 31432 20896
rect 31665 20893 31677 20896
rect 31711 20893 31723 20927
rect 31665 20887 31723 20893
rect 32493 20927 32551 20933
rect 32493 20893 32505 20927
rect 32539 20893 32551 20927
rect 32493 20887 32551 20893
rect 32508 20856 32536 20887
rect 32582 20884 32588 20936
rect 32640 20924 32646 20936
rect 32677 20927 32735 20933
rect 32677 20924 32689 20927
rect 32640 20896 32689 20924
rect 32640 20884 32646 20896
rect 32677 20893 32689 20896
rect 32723 20893 32735 20927
rect 32677 20887 32735 20893
rect 32766 20884 32772 20936
rect 32824 20924 32830 20936
rect 33612 20924 33640 20955
rect 34422 20952 34428 20964
rect 34480 20952 34486 21004
rect 34514 20952 34520 21004
rect 34572 20992 34578 21004
rect 34701 20995 34759 21001
rect 34701 20992 34713 20995
rect 34572 20964 34713 20992
rect 34572 20952 34578 20964
rect 34701 20961 34713 20964
rect 34747 20961 34759 20995
rect 34701 20955 34759 20961
rect 33778 20924 33784 20936
rect 32824 20896 33640 20924
rect 33739 20896 33784 20924
rect 32824 20884 32830 20896
rect 33778 20884 33784 20896
rect 33836 20884 33842 20936
rect 33965 20927 34023 20933
rect 33965 20893 33977 20927
rect 34011 20893 34023 20927
rect 33965 20887 34023 20893
rect 33042 20856 33048 20868
rect 32508 20828 33048 20856
rect 33042 20816 33048 20828
rect 33100 20816 33106 20868
rect 33980 20856 34008 20887
rect 34054 20884 34060 20936
rect 34112 20924 34118 20936
rect 34112 20896 34157 20924
rect 34112 20884 34118 20896
rect 34606 20884 34612 20936
rect 34664 20924 34670 20936
rect 35069 20927 35127 20933
rect 35069 20924 35081 20927
rect 34664 20896 35081 20924
rect 34664 20884 34670 20896
rect 35069 20893 35081 20896
rect 35115 20893 35127 20927
rect 35069 20887 35127 20893
rect 35161 20927 35219 20933
rect 35161 20893 35173 20927
rect 35207 20893 35219 20927
rect 35161 20887 35219 20893
rect 34790 20856 34796 20868
rect 33980 20828 34796 20856
rect 34790 20816 34796 20828
rect 34848 20816 34854 20868
rect 30892 20760 31432 20788
rect 30892 20748 30898 20760
rect 31846 20748 31852 20800
rect 31904 20788 31910 20800
rect 32309 20791 32367 20797
rect 32309 20788 32321 20791
rect 31904 20760 32321 20788
rect 31904 20748 31910 20760
rect 32309 20757 32321 20760
rect 32355 20757 32367 20791
rect 32309 20751 32367 20757
rect 33686 20748 33692 20800
rect 33744 20788 33750 20800
rect 35176 20788 35204 20887
rect 35866 20856 35894 21032
rect 38102 20992 38108 21004
rect 38063 20964 38108 20992
rect 38102 20952 38108 20964
rect 38160 20952 38166 21004
rect 36262 20924 36268 20936
rect 36223 20896 36268 20924
rect 36262 20884 36268 20896
rect 36320 20884 36326 20936
rect 36449 20859 36507 20865
rect 36449 20856 36461 20859
rect 35866 20828 36461 20856
rect 36449 20825 36461 20828
rect 36495 20825 36507 20859
rect 36449 20819 36507 20825
rect 35342 20788 35348 20800
rect 33744 20760 35204 20788
rect 35303 20760 35348 20788
rect 33744 20748 33750 20760
rect 35342 20748 35348 20760
rect 35400 20748 35406 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 2314 20544 2320 20596
rect 2372 20584 2378 20596
rect 26234 20584 26240 20596
rect 2372 20556 6914 20584
rect 2372 20544 2378 20556
rect 6886 20380 6914 20556
rect 12406 20556 26240 20584
rect 7834 20476 7840 20528
rect 7892 20516 7898 20528
rect 7929 20519 7987 20525
rect 7929 20516 7941 20519
rect 7892 20488 7941 20516
rect 7892 20476 7898 20488
rect 7929 20485 7941 20488
rect 7975 20485 7987 20519
rect 7929 20479 7987 20485
rect 9214 20380 9220 20392
rect 6886 20352 9220 20380
rect 9214 20340 9220 20352
rect 9272 20380 9278 20392
rect 9585 20383 9643 20389
rect 9585 20380 9597 20383
rect 9272 20352 9597 20380
rect 9272 20340 9278 20352
rect 9585 20349 9597 20352
rect 9631 20380 9643 20383
rect 12406 20380 12434 20556
rect 26234 20544 26240 20556
rect 26292 20544 26298 20596
rect 26418 20584 26424 20596
rect 26379 20556 26424 20584
rect 26418 20544 26424 20556
rect 26476 20544 26482 20596
rect 29549 20587 29607 20593
rect 29549 20553 29561 20587
rect 29595 20584 29607 20587
rect 29914 20584 29920 20596
rect 29595 20556 29920 20584
rect 29595 20553 29607 20556
rect 29549 20547 29607 20553
rect 29914 20544 29920 20556
rect 29972 20544 29978 20596
rect 30006 20544 30012 20596
rect 30064 20584 30070 20596
rect 33042 20584 33048 20596
rect 30064 20556 32904 20584
rect 33003 20556 33048 20584
rect 30064 20544 30070 20556
rect 15746 20516 15752 20528
rect 15659 20488 15752 20516
rect 15746 20476 15752 20488
rect 15804 20516 15810 20528
rect 16482 20516 16488 20528
rect 15804 20488 16488 20516
rect 15804 20476 15810 20488
rect 16482 20476 16488 20488
rect 16540 20476 16546 20528
rect 17773 20519 17831 20525
rect 17773 20516 17785 20519
rect 16868 20488 17785 20516
rect 15565 20451 15623 20457
rect 15565 20417 15577 20451
rect 15611 20448 15623 20451
rect 15654 20448 15660 20460
rect 15611 20420 15660 20448
rect 15611 20417 15623 20420
rect 15565 20411 15623 20417
rect 9631 20352 12434 20380
rect 9631 20349 9643 20352
rect 9585 20343 9643 20349
rect 15580 20312 15608 20411
rect 15654 20408 15660 20420
rect 15712 20408 15718 20460
rect 15838 20408 15844 20460
rect 15896 20448 15902 20460
rect 16868 20457 16896 20488
rect 17773 20485 17785 20488
rect 17819 20485 17831 20519
rect 17773 20479 17831 20485
rect 22094 20476 22100 20528
rect 22152 20516 22158 20528
rect 22830 20516 22836 20528
rect 22152 20488 22836 20516
rect 22152 20476 22158 20488
rect 22830 20476 22836 20488
rect 22888 20525 22894 20528
rect 22888 20519 22951 20525
rect 22888 20485 22905 20519
rect 22939 20516 22951 20519
rect 23109 20519 23167 20525
rect 22939 20485 22968 20516
rect 22888 20479 22968 20485
rect 23109 20485 23121 20519
rect 23155 20516 23167 20519
rect 23290 20516 23296 20528
rect 23155 20488 23296 20516
rect 23155 20485 23167 20488
rect 23109 20479 23167 20485
rect 22888 20476 22894 20479
rect 16669 20451 16727 20457
rect 16669 20448 16681 20451
rect 15896 20420 16681 20448
rect 15896 20408 15902 20420
rect 16669 20417 16681 20420
rect 16715 20417 16727 20451
rect 16669 20411 16727 20417
rect 16853 20451 16911 20457
rect 16853 20417 16865 20451
rect 16899 20417 16911 20451
rect 17494 20448 17500 20460
rect 17455 20420 17500 20448
rect 16853 20411 16911 20417
rect 17494 20408 17500 20420
rect 17552 20408 17558 20460
rect 17773 20383 17831 20389
rect 17773 20349 17785 20383
rect 17819 20380 17831 20383
rect 18598 20380 18604 20392
rect 17819 20352 18604 20380
rect 17819 20349 17831 20352
rect 17773 20343 17831 20349
rect 18598 20340 18604 20352
rect 18656 20340 18662 20392
rect 22940 20380 22968 20479
rect 23290 20476 23296 20488
rect 23348 20516 23354 20528
rect 23753 20519 23811 20525
rect 23753 20516 23765 20519
rect 23348 20488 23765 20516
rect 23348 20476 23354 20488
rect 23753 20485 23765 20488
rect 23799 20485 23811 20519
rect 23753 20479 23811 20485
rect 25308 20519 25366 20525
rect 25308 20485 25320 20519
rect 25354 20516 25366 20519
rect 27065 20519 27123 20525
rect 27065 20516 27077 20519
rect 25354 20488 27077 20516
rect 25354 20485 25366 20488
rect 25308 20479 25366 20485
rect 27065 20485 27077 20488
rect 27111 20485 27123 20519
rect 27065 20479 27123 20485
rect 29825 20519 29883 20525
rect 29825 20485 29837 20519
rect 29871 20516 29883 20519
rect 30024 20516 30052 20544
rect 29871 20488 30052 20516
rect 29871 20485 29883 20488
rect 29825 20479 29883 20485
rect 30374 20476 30380 20528
rect 30432 20516 30438 20528
rect 31662 20516 31668 20528
rect 30432 20488 31668 20516
rect 30432 20476 30438 20488
rect 31662 20476 31668 20488
rect 31720 20516 31726 20528
rect 32876 20516 32904 20556
rect 33042 20544 33048 20556
rect 33100 20544 33106 20596
rect 33686 20584 33692 20596
rect 33647 20556 33692 20584
rect 33686 20544 33692 20556
rect 33744 20544 33750 20596
rect 34054 20544 34060 20596
rect 34112 20584 34118 20596
rect 34241 20587 34299 20593
rect 34241 20584 34253 20587
rect 34112 20556 34253 20584
rect 34112 20544 34118 20556
rect 34241 20553 34253 20556
rect 34287 20553 34299 20587
rect 34241 20547 34299 20553
rect 33134 20516 33140 20528
rect 31720 20488 32720 20516
rect 32876 20488 33140 20516
rect 31720 20476 31726 20488
rect 23014 20408 23020 20460
rect 23072 20448 23078 20460
rect 23382 20448 23388 20460
rect 23072 20420 23388 20448
rect 23072 20408 23078 20420
rect 23382 20408 23388 20420
rect 23440 20448 23446 20460
rect 23569 20451 23627 20457
rect 23569 20448 23581 20451
rect 23440 20420 23581 20448
rect 23440 20408 23446 20420
rect 23569 20417 23581 20420
rect 23615 20417 23627 20451
rect 23569 20411 23627 20417
rect 23845 20451 23903 20457
rect 23845 20417 23857 20451
rect 23891 20417 23903 20451
rect 25038 20448 25044 20460
rect 24999 20420 25044 20448
rect 23845 20411 23903 20417
rect 23860 20380 23888 20411
rect 25038 20408 25044 20420
rect 25096 20408 25102 20460
rect 26970 20448 26976 20460
rect 26931 20420 26976 20448
rect 26970 20408 26976 20420
rect 27028 20408 27034 20460
rect 27154 20448 27160 20460
rect 27115 20420 27160 20448
rect 27154 20408 27160 20420
rect 27212 20408 27218 20460
rect 27890 20408 27896 20460
rect 27948 20448 27954 20460
rect 29730 20457 29736 20460
rect 28629 20451 28687 20457
rect 28629 20448 28641 20451
rect 27948 20420 28641 20448
rect 27948 20408 27954 20420
rect 28629 20417 28641 20420
rect 28675 20417 28687 20451
rect 28629 20411 28687 20417
rect 28721 20451 28779 20457
rect 28721 20417 28733 20451
rect 28767 20448 28779 20451
rect 29687 20451 29736 20457
rect 29687 20448 29699 20451
rect 28767 20420 29699 20448
rect 28767 20417 28779 20420
rect 28721 20411 28779 20417
rect 29687 20417 29699 20420
rect 29733 20417 29736 20451
rect 29687 20411 29736 20417
rect 29730 20408 29736 20411
rect 29788 20408 29794 20460
rect 29914 20408 29920 20460
rect 29972 20448 29978 20460
rect 30100 20451 30158 20457
rect 29972 20420 30017 20448
rect 29972 20408 29978 20420
rect 30100 20417 30112 20451
rect 30146 20417 30158 20451
rect 30100 20411 30158 20417
rect 22940 20352 23888 20380
rect 29546 20340 29552 20392
rect 29604 20380 29610 20392
rect 30116 20380 30144 20411
rect 30190 20408 30196 20460
rect 30248 20448 30254 20460
rect 30926 20448 30932 20460
rect 30248 20420 30293 20448
rect 30887 20420 30932 20448
rect 30248 20408 30254 20420
rect 30926 20408 30932 20420
rect 30984 20408 30990 20460
rect 32692 20457 32720 20488
rect 33134 20476 33140 20488
rect 33192 20476 33198 20528
rect 32677 20451 32735 20457
rect 32677 20417 32689 20451
rect 32723 20417 32735 20451
rect 32677 20411 32735 20417
rect 32861 20451 32919 20457
rect 32861 20417 32873 20451
rect 32907 20448 32919 20451
rect 33597 20451 33655 20457
rect 33597 20448 33609 20451
rect 32907 20420 33609 20448
rect 32907 20417 32919 20420
rect 32861 20411 32919 20417
rect 33597 20417 33609 20420
rect 33643 20448 33655 20451
rect 34330 20448 34336 20460
rect 33643 20420 34336 20448
rect 33643 20417 33655 20420
rect 33597 20411 33655 20417
rect 34330 20408 34336 20420
rect 34388 20448 34394 20460
rect 34425 20451 34483 20457
rect 34425 20448 34437 20451
rect 34388 20420 34437 20448
rect 34388 20408 34394 20420
rect 34425 20417 34437 20420
rect 34471 20448 34483 20451
rect 35526 20448 35532 20460
rect 34471 20420 35532 20448
rect 34471 20417 34483 20420
rect 34425 20411 34483 20417
rect 35526 20408 35532 20420
rect 35584 20408 35590 20460
rect 36262 20408 36268 20460
rect 36320 20448 36326 20460
rect 36541 20451 36599 20457
rect 36541 20448 36553 20451
rect 36320 20420 36553 20448
rect 36320 20408 36326 20420
rect 36541 20417 36553 20420
rect 36587 20417 36599 20451
rect 36541 20411 36599 20417
rect 37369 20451 37427 20457
rect 37369 20417 37381 20451
rect 37415 20448 37427 20451
rect 38194 20448 38200 20460
rect 37415 20420 38200 20448
rect 37415 20417 37427 20420
rect 37369 20411 37427 20417
rect 38194 20408 38200 20420
rect 38252 20408 38258 20460
rect 29604 20352 30144 20380
rect 31021 20383 31079 20389
rect 29604 20340 29610 20352
rect 31021 20349 31033 20383
rect 31067 20380 31079 20383
rect 31067 20352 33088 20380
rect 31067 20349 31079 20352
rect 31021 20343 31079 20349
rect 23014 20312 23020 20324
rect 15580 20284 23020 20312
rect 23014 20272 23020 20284
rect 23072 20272 23078 20324
rect 31297 20315 31355 20321
rect 31297 20281 31309 20315
rect 31343 20312 31355 20315
rect 31754 20312 31760 20324
rect 31343 20284 31760 20312
rect 31343 20281 31355 20284
rect 31297 20275 31355 20281
rect 31754 20272 31760 20284
rect 31812 20272 31818 20324
rect 33060 20312 33088 20352
rect 33134 20340 33140 20392
rect 33192 20380 33198 20392
rect 34701 20383 34759 20389
rect 34701 20380 34713 20383
rect 33192 20352 34713 20380
rect 33192 20340 33198 20352
rect 34701 20349 34713 20352
rect 34747 20349 34759 20383
rect 34701 20343 34759 20349
rect 33686 20312 33692 20324
rect 33060 20284 33692 20312
rect 33686 20272 33692 20284
rect 33744 20272 33750 20324
rect 34606 20312 34612 20324
rect 34567 20284 34612 20312
rect 34606 20272 34612 20284
rect 34664 20272 34670 20324
rect 1394 20204 1400 20256
rect 1452 20244 1458 20256
rect 1581 20247 1639 20253
rect 1581 20244 1593 20247
rect 1452 20216 1593 20244
rect 1452 20204 1458 20216
rect 1581 20213 1593 20216
rect 1627 20213 1639 20247
rect 1581 20207 1639 20213
rect 15470 20204 15476 20256
rect 15528 20244 15534 20256
rect 15565 20247 15623 20253
rect 15565 20244 15577 20247
rect 15528 20216 15577 20244
rect 15528 20204 15534 20216
rect 15565 20213 15577 20216
rect 15611 20213 15623 20247
rect 16850 20244 16856 20256
rect 16811 20216 16856 20244
rect 15565 20207 15623 20213
rect 16850 20204 16856 20216
rect 16908 20204 16914 20256
rect 17589 20247 17647 20253
rect 17589 20213 17601 20247
rect 17635 20244 17647 20247
rect 17954 20244 17960 20256
rect 17635 20216 17960 20244
rect 17635 20213 17647 20216
rect 17589 20207 17647 20213
rect 17954 20204 17960 20216
rect 18012 20204 18018 20256
rect 21818 20204 21824 20256
rect 21876 20244 21882 20256
rect 22741 20247 22799 20253
rect 22741 20244 22753 20247
rect 21876 20216 22753 20244
rect 21876 20204 21882 20216
rect 22741 20213 22753 20216
rect 22787 20213 22799 20247
rect 22922 20244 22928 20256
rect 22883 20216 22928 20244
rect 22741 20207 22799 20213
rect 22922 20204 22928 20216
rect 22980 20204 22986 20256
rect 23566 20244 23572 20256
rect 23527 20216 23572 20244
rect 23566 20204 23572 20216
rect 23624 20204 23630 20256
rect 26234 20204 26240 20256
rect 26292 20244 26298 20256
rect 32490 20244 32496 20256
rect 26292 20216 32496 20244
rect 26292 20204 26298 20216
rect 32490 20204 32496 20216
rect 32548 20204 32554 20256
rect 37461 20247 37519 20253
rect 37461 20213 37473 20247
rect 37507 20244 37519 20247
rect 37918 20244 37924 20256
rect 37507 20216 37924 20244
rect 37507 20213 37519 20216
rect 37461 20207 37519 20213
rect 37918 20204 37924 20216
rect 37976 20204 37982 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 15565 20043 15623 20049
rect 15565 20009 15577 20043
rect 15611 20040 15623 20043
rect 15746 20040 15752 20052
rect 15611 20012 15752 20040
rect 15611 20009 15623 20012
rect 15565 20003 15623 20009
rect 15746 20000 15752 20012
rect 15804 20000 15810 20052
rect 15838 20000 15844 20052
rect 15896 20040 15902 20052
rect 17865 20043 17923 20049
rect 17865 20040 17877 20043
rect 15896 20012 17877 20040
rect 15896 20000 15902 20012
rect 17865 20009 17877 20012
rect 17911 20009 17923 20043
rect 18046 20040 18052 20052
rect 18007 20012 18052 20040
rect 17865 20003 17923 20009
rect 18046 20000 18052 20012
rect 18104 20000 18110 20052
rect 19705 20043 19763 20049
rect 19705 20009 19717 20043
rect 19751 20040 19763 20043
rect 20346 20040 20352 20052
rect 19751 20012 20352 20040
rect 19751 20009 19763 20012
rect 19705 20003 19763 20009
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 29733 20043 29791 20049
rect 29733 20009 29745 20043
rect 29779 20040 29791 20043
rect 30282 20040 30288 20052
rect 29779 20012 30288 20040
rect 29779 20009 29791 20012
rect 29733 20003 29791 20009
rect 30282 20000 30288 20012
rect 30340 20000 30346 20052
rect 30745 20043 30803 20049
rect 30745 20009 30757 20043
rect 30791 20040 30803 20043
rect 30926 20040 30932 20052
rect 30791 20012 30932 20040
rect 30791 20009 30803 20012
rect 30745 20003 30803 20009
rect 30926 20000 30932 20012
rect 30984 20000 30990 20052
rect 32401 20043 32459 20049
rect 32401 20009 32413 20043
rect 32447 20040 32459 20043
rect 33318 20040 33324 20052
rect 32447 20012 33324 20040
rect 32447 20009 32459 20012
rect 32401 20003 32459 20009
rect 33318 20000 33324 20012
rect 33376 20000 33382 20052
rect 21913 19975 21971 19981
rect 21913 19941 21925 19975
rect 21959 19972 21971 19975
rect 23566 19972 23572 19984
rect 21959 19944 23572 19972
rect 21959 19941 21971 19944
rect 21913 19935 21971 19941
rect 23566 19932 23572 19944
rect 23624 19932 23630 19984
rect 1394 19904 1400 19916
rect 1355 19876 1400 19904
rect 1394 19864 1400 19876
rect 1452 19864 1458 19916
rect 1854 19904 1860 19916
rect 1815 19876 1860 19904
rect 1854 19864 1860 19876
rect 1912 19864 1918 19916
rect 14182 19904 14188 19916
rect 14143 19876 14188 19904
rect 14182 19864 14188 19876
rect 14240 19864 14246 19916
rect 18598 19864 18604 19916
rect 18656 19904 18662 19916
rect 20162 19904 20168 19916
rect 18656 19876 20168 19904
rect 18656 19864 18662 19876
rect 20162 19864 20168 19876
rect 20220 19904 20226 19916
rect 20625 19907 20683 19913
rect 20625 19904 20637 19907
rect 20220 19876 20637 19904
rect 20220 19864 20226 19876
rect 20625 19873 20637 19876
rect 20671 19873 20683 19907
rect 20625 19867 20683 19873
rect 22370 19864 22376 19916
rect 22428 19904 22434 19916
rect 22557 19907 22615 19913
rect 22557 19904 22569 19907
rect 22428 19876 22569 19904
rect 22428 19864 22434 19876
rect 22557 19873 22569 19876
rect 22603 19873 22615 19907
rect 22830 19904 22836 19916
rect 22791 19876 22836 19904
rect 22557 19867 22615 19873
rect 22830 19864 22836 19876
rect 22888 19864 22894 19916
rect 26694 19864 26700 19916
rect 26752 19904 26758 19916
rect 27341 19907 27399 19913
rect 27341 19904 27353 19907
rect 26752 19876 27353 19904
rect 26752 19864 26758 19876
rect 27341 19873 27353 19876
rect 27387 19873 27399 19907
rect 37182 19904 37188 19916
rect 37143 19876 37188 19904
rect 27341 19867 27399 19873
rect 37182 19864 37188 19876
rect 37240 19864 37246 19916
rect 37918 19904 37924 19916
rect 37879 19876 37924 19904
rect 37918 19864 37924 19876
rect 37976 19864 37982 19916
rect 7745 19839 7803 19845
rect 7745 19805 7757 19839
rect 7791 19836 7803 19839
rect 7834 19836 7840 19848
rect 7791 19808 7840 19836
rect 7791 19805 7803 19808
rect 7745 19799 7803 19805
rect 7834 19796 7840 19808
rect 7892 19796 7898 19848
rect 14200 19836 14228 19864
rect 16025 19839 16083 19845
rect 16025 19836 16037 19839
rect 14200 19808 16037 19836
rect 16025 19805 16037 19808
rect 16071 19836 16083 19839
rect 17034 19836 17040 19848
rect 16071 19808 17040 19836
rect 16071 19805 16083 19808
rect 16025 19799 16083 19805
rect 17034 19796 17040 19808
rect 17092 19836 17098 19848
rect 17862 19836 17868 19848
rect 17092 19808 17868 19836
rect 17092 19796 17098 19808
rect 17862 19796 17868 19808
rect 17920 19796 17926 19848
rect 20346 19836 20352 19848
rect 20307 19808 20352 19836
rect 20346 19796 20352 19808
rect 20404 19796 20410 19848
rect 20441 19839 20499 19845
rect 20441 19805 20453 19839
rect 20487 19836 20499 19839
rect 21818 19836 21824 19848
rect 20487 19808 21824 19836
rect 20487 19805 20499 19808
rect 20441 19799 20499 19805
rect 1581 19771 1639 19777
rect 1581 19737 1593 19771
rect 1627 19768 1639 19771
rect 1946 19768 1952 19780
rect 1627 19740 1952 19768
rect 1627 19737 1639 19740
rect 1581 19731 1639 19737
rect 1946 19728 1952 19740
rect 2004 19728 2010 19780
rect 8110 19768 8116 19780
rect 8071 19740 8116 19768
rect 8110 19728 8116 19740
rect 8168 19728 8174 19780
rect 14452 19771 14510 19777
rect 14452 19737 14464 19771
rect 14498 19768 14510 19771
rect 15286 19768 15292 19780
rect 14498 19740 15292 19768
rect 14498 19737 14510 19740
rect 14452 19731 14510 19737
rect 15286 19728 15292 19740
rect 15344 19728 15350 19780
rect 16292 19771 16350 19777
rect 16292 19737 16304 19771
rect 16338 19768 16350 19771
rect 16850 19768 16856 19780
rect 16338 19740 16856 19768
rect 16338 19737 16350 19740
rect 16292 19731 16350 19737
rect 16850 19728 16856 19740
rect 16908 19728 16914 19780
rect 17494 19768 17500 19780
rect 17407 19740 17500 19768
rect 17420 19709 17448 19740
rect 17494 19728 17500 19740
rect 17552 19768 17558 19780
rect 18233 19771 18291 19777
rect 18233 19768 18245 19771
rect 17552 19740 18245 19768
rect 17552 19728 17558 19740
rect 18233 19737 18245 19740
rect 18279 19737 18291 19771
rect 18233 19731 18291 19737
rect 19426 19728 19432 19780
rect 19484 19768 19490 19780
rect 19889 19771 19947 19777
rect 19889 19768 19901 19771
rect 19484 19740 19901 19768
rect 19484 19728 19490 19740
rect 19889 19737 19901 19740
rect 19935 19737 19947 19771
rect 19889 19731 19947 19737
rect 17405 19703 17463 19709
rect 17405 19669 17417 19703
rect 17451 19669 17463 19703
rect 17405 19663 17463 19669
rect 18033 19703 18091 19709
rect 18033 19669 18045 19703
rect 18079 19700 18091 19703
rect 19242 19700 19248 19712
rect 18079 19672 19248 19700
rect 18079 19669 18091 19672
rect 18033 19663 18091 19669
rect 19242 19660 19248 19672
rect 19300 19700 19306 19712
rect 19521 19703 19579 19709
rect 19521 19700 19533 19703
rect 19300 19672 19533 19700
rect 19300 19660 19306 19672
rect 19521 19669 19533 19672
rect 19567 19669 19579 19703
rect 19521 19663 19579 19669
rect 19689 19703 19747 19709
rect 19689 19669 19701 19703
rect 19735 19700 19747 19703
rect 20070 19700 20076 19712
rect 19735 19672 20076 19700
rect 19735 19669 19747 19672
rect 19689 19663 19747 19669
rect 20070 19660 20076 19672
rect 20128 19700 20134 19712
rect 20456 19700 20484 19799
rect 21818 19796 21824 19808
rect 21876 19796 21882 19848
rect 22097 19839 22155 19845
rect 22097 19805 22109 19839
rect 22143 19836 22155 19839
rect 24946 19836 24952 19848
rect 22143 19808 24952 19836
rect 22143 19805 22155 19808
rect 22097 19799 22155 19805
rect 24946 19796 24952 19808
rect 25004 19836 25010 19848
rect 25041 19839 25099 19845
rect 25041 19836 25053 19839
rect 25004 19808 25053 19836
rect 25004 19796 25010 19808
rect 25041 19805 25053 19808
rect 25087 19805 25099 19839
rect 25041 19799 25099 19805
rect 26970 19796 26976 19848
rect 27028 19836 27034 19848
rect 27525 19839 27583 19845
rect 27525 19836 27537 19839
rect 27028 19808 27537 19836
rect 27028 19796 27034 19808
rect 27525 19805 27537 19808
rect 27571 19805 27583 19839
rect 27525 19799 27583 19805
rect 27614 19796 27620 19848
rect 27672 19836 27678 19848
rect 28077 19839 28135 19845
rect 27672 19808 27717 19836
rect 27672 19796 27678 19808
rect 28077 19805 28089 19839
rect 28123 19805 28135 19839
rect 28077 19799 28135 19805
rect 24854 19768 24860 19780
rect 24815 19740 24860 19768
rect 24854 19728 24860 19740
rect 24912 19768 24918 19780
rect 27341 19771 27399 19777
rect 24912 19740 27108 19768
rect 24912 19728 24918 19740
rect 20128 19672 20484 19700
rect 20625 19703 20683 19709
rect 20128 19660 20134 19672
rect 20625 19669 20637 19703
rect 20671 19700 20683 19703
rect 20898 19700 20904 19712
rect 20671 19672 20904 19700
rect 20671 19669 20683 19672
rect 20625 19663 20683 19669
rect 20898 19660 20904 19672
rect 20956 19660 20962 19712
rect 21821 19703 21879 19709
rect 21821 19669 21833 19703
rect 21867 19700 21879 19703
rect 24762 19700 24768 19712
rect 21867 19672 24768 19700
rect 21867 19669 21879 19672
rect 21821 19663 21879 19669
rect 24762 19660 24768 19672
rect 24820 19660 24826 19712
rect 26142 19660 26148 19712
rect 26200 19700 26206 19712
rect 26252 19700 26280 19740
rect 26200 19672 26280 19700
rect 27080 19700 27108 19740
rect 27341 19737 27353 19771
rect 27387 19768 27399 19771
rect 28092 19768 28120 19799
rect 28166 19796 28172 19848
rect 28224 19836 28230 19848
rect 28261 19839 28319 19845
rect 28261 19836 28273 19839
rect 28224 19808 28273 19836
rect 28224 19796 28230 19808
rect 28261 19805 28273 19808
rect 28307 19805 28319 19839
rect 28261 19799 28319 19805
rect 28902 19796 28908 19848
rect 28960 19836 28966 19848
rect 29641 19839 29699 19845
rect 29641 19836 29653 19839
rect 28960 19808 29653 19836
rect 28960 19796 28966 19808
rect 29641 19805 29653 19808
rect 29687 19805 29699 19839
rect 30834 19836 30840 19848
rect 30795 19808 30840 19836
rect 29641 19799 29699 19805
rect 30834 19796 30840 19808
rect 30892 19796 30898 19848
rect 31662 19796 31668 19848
rect 31720 19836 31726 19848
rect 32217 19839 32275 19845
rect 32217 19836 32229 19839
rect 31720 19808 32229 19836
rect 31720 19796 31726 19808
rect 32217 19805 32229 19808
rect 32263 19805 32275 19839
rect 32217 19799 32275 19805
rect 32401 19839 32459 19845
rect 32401 19805 32413 19839
rect 32447 19836 32459 19839
rect 33686 19836 33692 19848
rect 32447 19808 33692 19836
rect 32447 19805 32459 19808
rect 32401 19799 32459 19805
rect 33686 19796 33692 19808
rect 33744 19796 33750 19848
rect 38102 19796 38108 19848
rect 38160 19836 38166 19848
rect 38160 19808 38205 19836
rect 38160 19796 38166 19808
rect 27387 19740 28120 19768
rect 27387 19737 27399 19740
rect 27341 19731 27399 19737
rect 27798 19700 27804 19712
rect 27080 19672 27804 19700
rect 26200 19660 26206 19672
rect 27798 19660 27804 19672
rect 27856 19660 27862 19712
rect 28169 19703 28227 19709
rect 28169 19669 28181 19703
rect 28215 19700 28227 19703
rect 28258 19700 28264 19712
rect 28215 19672 28264 19700
rect 28215 19669 28227 19672
rect 28169 19663 28227 19669
rect 28258 19660 28264 19672
rect 28316 19660 28322 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 16758 19496 16764 19508
rect 6886 19468 16764 19496
rect 2038 19360 2044 19372
rect 1951 19332 2044 19360
rect 2038 19320 2044 19332
rect 2096 19360 2102 19372
rect 6886 19360 6914 19468
rect 16758 19456 16764 19468
rect 16816 19456 16822 19508
rect 17589 19499 17647 19505
rect 17589 19465 17601 19499
rect 17635 19496 17647 19499
rect 17954 19496 17960 19508
rect 17635 19468 17960 19496
rect 17635 19465 17647 19468
rect 17589 19459 17647 19465
rect 17954 19456 17960 19468
rect 18012 19456 18018 19508
rect 18049 19499 18107 19505
rect 18049 19465 18061 19499
rect 18095 19496 18107 19499
rect 19426 19496 19432 19508
rect 18095 19468 19432 19496
rect 18095 19465 18107 19468
rect 18049 19459 18107 19465
rect 19426 19456 19432 19468
rect 19484 19456 19490 19508
rect 19889 19499 19947 19505
rect 19889 19465 19901 19499
rect 19935 19496 19947 19499
rect 20346 19496 20352 19508
rect 19935 19468 20352 19496
rect 19935 19465 19947 19468
rect 19889 19459 19947 19465
rect 20346 19456 20352 19468
rect 20404 19456 20410 19508
rect 22370 19456 22376 19508
rect 22428 19496 22434 19508
rect 23201 19499 23259 19505
rect 23201 19496 23213 19499
rect 22428 19468 23213 19496
rect 22428 19456 22434 19468
rect 23201 19465 23213 19468
rect 23247 19465 23259 19499
rect 23201 19459 23259 19465
rect 23382 19456 23388 19508
rect 23440 19496 23446 19508
rect 23661 19499 23719 19505
rect 23661 19496 23673 19499
rect 23440 19468 23673 19496
rect 23440 19456 23446 19468
rect 23661 19465 23673 19468
rect 23707 19465 23719 19499
rect 26970 19496 26976 19508
rect 26931 19468 26976 19496
rect 23661 19459 23719 19465
rect 26970 19456 26976 19468
rect 27028 19456 27034 19508
rect 27614 19456 27620 19508
rect 27672 19496 27678 19508
rect 28902 19496 28908 19508
rect 27672 19468 28908 19496
rect 27672 19456 27678 19468
rect 28902 19456 28908 19468
rect 28960 19496 28966 19508
rect 29365 19499 29423 19505
rect 29365 19496 29377 19499
rect 28960 19468 29377 19496
rect 28960 19456 28966 19468
rect 29365 19465 29377 19468
rect 29411 19465 29423 19499
rect 29365 19459 29423 19465
rect 17862 19388 17868 19440
rect 17920 19428 17926 19440
rect 22278 19428 22284 19440
rect 17920 19400 21312 19428
rect 17920 19388 17926 19400
rect 15470 19360 15476 19372
rect 2096 19332 6914 19360
rect 15431 19332 15476 19360
rect 2096 19320 2102 19332
rect 15470 19320 15476 19332
rect 15528 19320 15534 19372
rect 15657 19363 15715 19369
rect 15657 19329 15669 19363
rect 15703 19360 15715 19363
rect 15838 19360 15844 19372
rect 15703 19332 15844 19360
rect 15703 19329 15715 19332
rect 15657 19323 15715 19329
rect 15838 19320 15844 19332
rect 15896 19320 15902 19372
rect 17405 19363 17463 19369
rect 17405 19329 17417 19363
rect 17451 19360 17463 19363
rect 17954 19360 17960 19372
rect 17451 19332 17960 19360
rect 17451 19329 17463 19332
rect 17405 19323 17463 19329
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 19173 19363 19231 19369
rect 19173 19329 19185 19363
rect 19219 19360 19231 19363
rect 19334 19360 19340 19372
rect 19219 19332 19340 19360
rect 19219 19329 19231 19332
rect 19173 19323 19231 19329
rect 19334 19320 19340 19332
rect 19392 19320 19398 19372
rect 19444 19369 19472 19400
rect 19429 19363 19487 19369
rect 19429 19329 19441 19363
rect 19475 19329 19487 19363
rect 20990 19360 20996 19372
rect 21048 19369 21054 19372
rect 21284 19369 21312 19400
rect 21836 19400 22284 19428
rect 21836 19369 21864 19400
rect 22278 19388 22284 19400
rect 22336 19388 22342 19440
rect 24762 19388 24768 19440
rect 24820 19437 24826 19440
rect 24820 19428 24832 19437
rect 24820 19400 24865 19428
rect 24820 19391 24832 19400
rect 24820 19388 24826 19391
rect 22094 19369 22100 19372
rect 20960 19332 20996 19360
rect 19429 19323 19487 19329
rect 20990 19320 20996 19332
rect 21048 19323 21060 19369
rect 21269 19363 21327 19369
rect 21269 19329 21281 19363
rect 21315 19360 21327 19363
rect 21821 19363 21879 19369
rect 21821 19360 21833 19363
rect 21315 19332 21833 19360
rect 21315 19329 21327 19332
rect 21269 19323 21327 19329
rect 21821 19329 21833 19332
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 22088 19323 22100 19369
rect 22152 19360 22158 19372
rect 25038 19360 25044 19372
rect 22152 19332 22188 19360
rect 24999 19332 25044 19360
rect 21048 19320 21054 19323
rect 22094 19320 22100 19323
rect 22152 19320 22158 19332
rect 25038 19320 25044 19332
rect 25096 19320 25102 19372
rect 26142 19320 26148 19372
rect 26200 19360 26206 19372
rect 26237 19363 26295 19369
rect 26237 19360 26249 19363
rect 26200 19332 26249 19360
rect 26200 19320 26206 19332
rect 26237 19329 26249 19332
rect 26283 19329 26295 19363
rect 26237 19323 26295 19329
rect 26421 19363 26479 19369
rect 26421 19329 26433 19363
rect 26467 19360 26479 19363
rect 26988 19360 27016 19456
rect 28534 19428 28540 19440
rect 28000 19400 28540 19428
rect 27154 19360 27160 19372
rect 26467 19332 27016 19360
rect 27115 19332 27160 19360
rect 26467 19329 26479 19332
rect 26421 19323 26479 19329
rect 27154 19320 27160 19332
rect 27212 19320 27218 19372
rect 28000 19369 28028 19400
rect 28534 19388 28540 19400
rect 28592 19388 28598 19440
rect 28258 19369 28264 19372
rect 27985 19363 28043 19369
rect 27985 19329 27997 19363
rect 28031 19329 28043 19363
rect 28252 19360 28264 19369
rect 28219 19332 28264 19360
rect 27985 19323 28043 19329
rect 28252 19323 28264 19332
rect 28258 19320 28264 19323
rect 28316 19320 28322 19372
rect 33134 19320 33140 19372
rect 33192 19360 33198 19372
rect 34238 19360 34244 19372
rect 33192 19332 34244 19360
rect 33192 19320 33198 19332
rect 34238 19320 34244 19332
rect 34296 19360 34302 19372
rect 34425 19363 34483 19369
rect 34425 19360 34437 19363
rect 34296 19332 34437 19360
rect 34296 19320 34302 19332
rect 34425 19329 34437 19332
rect 34471 19329 34483 19363
rect 34425 19323 34483 19329
rect 37829 19363 37887 19369
rect 37829 19329 37841 19363
rect 37875 19360 37887 19363
rect 38102 19360 38108 19372
rect 37875 19332 38108 19360
rect 37875 19329 37887 19332
rect 37829 19323 37887 19329
rect 38102 19320 38108 19332
rect 38160 19320 38166 19372
rect 15286 19292 15292 19304
rect 15247 19264 15292 19292
rect 15286 19252 15292 19264
rect 15344 19252 15350 19304
rect 15746 19292 15752 19304
rect 15707 19264 15752 19292
rect 15746 19252 15752 19264
rect 15804 19252 15810 19304
rect 17221 19295 17279 19301
rect 17221 19261 17233 19295
rect 17267 19292 17279 19295
rect 18138 19292 18144 19304
rect 17267 19264 18144 19292
rect 17267 19261 17279 19264
rect 17221 19255 17279 19261
rect 18138 19252 18144 19264
rect 18196 19252 18202 19304
rect 27341 19295 27399 19301
rect 27341 19261 27353 19295
rect 27387 19292 27399 19295
rect 27890 19292 27896 19304
rect 27387 19264 27896 19292
rect 27387 19261 27399 19264
rect 27341 19255 27399 19261
rect 27890 19252 27896 19264
rect 27948 19252 27954 19304
rect 33778 19252 33784 19304
rect 33836 19292 33842 19304
rect 34057 19295 34115 19301
rect 34057 19292 34069 19295
rect 33836 19264 34069 19292
rect 33836 19252 33842 19264
rect 34057 19261 34069 19264
rect 34103 19261 34115 19295
rect 34330 19292 34336 19304
rect 34291 19264 34336 19292
rect 34057 19255 34115 19261
rect 34330 19252 34336 19264
rect 34388 19252 34394 19304
rect 26421 19159 26479 19165
rect 26421 19125 26433 19159
rect 26467 19156 26479 19159
rect 26602 19156 26608 19168
rect 26467 19128 26608 19156
rect 26467 19125 26479 19128
rect 26421 19119 26479 19125
rect 26602 19116 26608 19128
rect 26660 19116 26666 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 17865 18955 17923 18961
rect 17865 18921 17877 18955
rect 17911 18952 17923 18955
rect 17954 18952 17960 18964
rect 17911 18924 17960 18952
rect 17911 18921 17923 18924
rect 17865 18915 17923 18921
rect 17954 18912 17960 18924
rect 18012 18952 18018 18964
rect 19242 18952 19248 18964
rect 18012 18924 19248 18952
rect 18012 18912 18018 18924
rect 19242 18912 19248 18924
rect 19300 18912 19306 18964
rect 19334 18912 19340 18964
rect 19392 18952 19398 18964
rect 19429 18955 19487 18961
rect 19429 18952 19441 18955
rect 19392 18924 19441 18952
rect 19392 18912 19398 18924
rect 19429 18921 19441 18924
rect 19475 18921 19487 18955
rect 19429 18915 19487 18921
rect 20901 18955 20959 18961
rect 20901 18921 20913 18955
rect 20947 18952 20959 18955
rect 20990 18952 20996 18964
rect 20947 18924 20996 18952
rect 20947 18921 20959 18924
rect 20901 18915 20959 18921
rect 20990 18912 20996 18924
rect 21048 18912 21054 18964
rect 22094 18952 22100 18964
rect 22055 18924 22100 18952
rect 22094 18912 22100 18924
rect 22152 18912 22158 18964
rect 22465 18955 22523 18961
rect 22465 18921 22477 18955
rect 22511 18952 22523 18955
rect 22830 18952 22836 18964
rect 22511 18924 22836 18952
rect 22511 18921 22523 18924
rect 22465 18915 22523 18921
rect 22830 18912 22836 18924
rect 22888 18912 22894 18964
rect 24854 18952 24860 18964
rect 22940 18924 24860 18952
rect 22940 18884 22968 18924
rect 24854 18912 24860 18924
rect 24912 18912 24918 18964
rect 27890 18952 27896 18964
rect 27851 18924 27896 18952
rect 27890 18912 27896 18924
rect 27948 18912 27954 18964
rect 28077 18955 28135 18961
rect 28077 18921 28089 18955
rect 28123 18952 28135 18955
rect 28166 18952 28172 18964
rect 28123 18924 28172 18952
rect 28123 18921 28135 18924
rect 28077 18915 28135 18921
rect 28166 18912 28172 18924
rect 28224 18952 28230 18964
rect 28905 18955 28963 18961
rect 28905 18952 28917 18955
rect 28224 18924 28917 18952
rect 28224 18912 28230 18924
rect 28905 18921 28917 18924
rect 28951 18952 28963 18955
rect 28951 18924 29868 18952
rect 28951 18921 28963 18924
rect 28905 18915 28963 18921
rect 18616 18856 22968 18884
rect 23017 18887 23075 18893
rect 17957 18819 18015 18825
rect 17957 18785 17969 18819
rect 18003 18816 18015 18819
rect 18138 18816 18144 18828
rect 18003 18788 18144 18816
rect 18003 18785 18015 18788
rect 17957 18779 18015 18785
rect 18138 18776 18144 18788
rect 18196 18776 18202 18828
rect 17681 18751 17739 18757
rect 17681 18717 17693 18751
rect 17727 18717 17739 18751
rect 17681 18711 17739 18717
rect 17696 18680 17724 18711
rect 18046 18708 18052 18760
rect 18104 18748 18110 18760
rect 18616 18757 18644 18856
rect 23017 18853 23029 18887
rect 23063 18853 23075 18887
rect 23017 18847 23075 18853
rect 20257 18819 20315 18825
rect 20257 18785 20269 18819
rect 20303 18816 20315 18819
rect 20346 18816 20352 18828
rect 20303 18788 20352 18816
rect 20303 18785 20315 18788
rect 20257 18779 20315 18785
rect 20346 18776 20352 18788
rect 20404 18776 20410 18828
rect 23032 18816 23060 18847
rect 22296 18788 23060 18816
rect 26881 18819 26939 18825
rect 18417 18751 18475 18757
rect 18417 18748 18429 18751
rect 18104 18720 18429 18748
rect 18104 18708 18110 18720
rect 18417 18717 18429 18720
rect 18463 18717 18475 18751
rect 18417 18711 18475 18717
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18717 18659 18751
rect 19242 18748 19248 18760
rect 19203 18720 19248 18748
rect 18601 18711 18659 18717
rect 19242 18708 19248 18720
rect 19300 18708 19306 18760
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 19392 18720 19441 18748
rect 19392 18708 19398 18720
rect 19429 18717 19441 18720
rect 19475 18717 19487 18751
rect 20070 18748 20076 18760
rect 20031 18720 20076 18748
rect 19429 18711 19487 18717
rect 20070 18708 20076 18720
rect 20128 18708 20134 18760
rect 20717 18751 20775 18757
rect 20717 18717 20729 18751
rect 20763 18717 20775 18751
rect 20898 18748 20904 18760
rect 20859 18720 20904 18748
rect 20717 18711 20775 18717
rect 18509 18683 18567 18689
rect 18509 18680 18521 18683
rect 17696 18652 18521 18680
rect 18509 18649 18521 18652
rect 18555 18649 18567 18683
rect 18509 18643 18567 18649
rect 19889 18683 19947 18689
rect 19889 18649 19901 18683
rect 19935 18680 19947 18683
rect 19978 18680 19984 18692
rect 19935 18652 19984 18680
rect 19935 18649 19947 18652
rect 19889 18643 19947 18649
rect 19978 18640 19984 18652
rect 20036 18680 20042 18692
rect 20732 18680 20760 18711
rect 20898 18708 20904 18720
rect 20956 18708 20962 18760
rect 22296 18757 22324 18788
rect 26881 18785 26893 18819
rect 26927 18816 26939 18819
rect 27246 18816 27252 18828
rect 26927 18788 27252 18816
rect 26927 18785 26939 18788
rect 26881 18779 26939 18785
rect 27246 18776 27252 18788
rect 27304 18816 27310 18828
rect 27908 18816 27936 18912
rect 29549 18887 29607 18893
rect 29549 18853 29561 18887
rect 29595 18853 29607 18887
rect 29549 18847 29607 18853
rect 29564 18816 29592 18847
rect 27304 18788 27936 18816
rect 28736 18788 29592 18816
rect 27304 18776 27310 18788
rect 22281 18751 22339 18757
rect 22281 18717 22293 18751
rect 22327 18717 22339 18751
rect 22281 18711 22339 18717
rect 22557 18751 22615 18757
rect 22557 18717 22569 18751
rect 22603 18717 22615 18751
rect 22557 18711 22615 18717
rect 20036 18652 20760 18680
rect 20036 18640 20042 18652
rect 17310 18572 17316 18624
rect 17368 18612 17374 18624
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 17368 18584 17509 18612
rect 17368 18572 17374 18584
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 22572 18612 22600 18711
rect 22830 18708 22836 18760
rect 22888 18748 22894 18760
rect 23293 18751 23351 18757
rect 23293 18748 23305 18751
rect 22888 18720 23305 18748
rect 22888 18708 22894 18720
rect 23293 18717 23305 18720
rect 23339 18717 23351 18751
rect 26602 18748 26608 18760
rect 26563 18720 26608 18748
rect 23293 18711 23351 18717
rect 26602 18708 26608 18720
rect 26660 18708 26666 18760
rect 26786 18748 26792 18760
rect 26747 18720 26792 18748
rect 26786 18708 26792 18720
rect 26844 18708 26850 18760
rect 28736 18757 28764 18788
rect 29840 18757 29868 18924
rect 31754 18816 31760 18828
rect 31715 18788 31760 18816
rect 31754 18776 31760 18788
rect 31812 18776 31818 18828
rect 33134 18816 33140 18828
rect 32876 18788 33140 18816
rect 28721 18751 28779 18757
rect 27540 18720 28212 18748
rect 23014 18680 23020 18692
rect 22975 18652 23020 18680
rect 23014 18640 23020 18652
rect 23072 18680 23078 18692
rect 27540 18680 27568 18720
rect 23072 18652 27568 18680
rect 23072 18640 23078 18652
rect 27614 18640 27620 18692
rect 27672 18680 27678 18692
rect 27709 18683 27767 18689
rect 27709 18680 27721 18683
rect 27672 18652 27721 18680
rect 27672 18640 27678 18652
rect 27709 18649 27721 18652
rect 27755 18649 27767 18683
rect 28184 18680 28212 18720
rect 28721 18717 28733 18751
rect 28767 18717 28779 18751
rect 28721 18711 28779 18717
rect 28997 18751 29055 18757
rect 28997 18717 29009 18751
rect 29043 18748 29055 18751
rect 29825 18751 29883 18757
rect 29043 18720 29776 18748
rect 29043 18717 29055 18720
rect 28997 18711 29055 18717
rect 29086 18680 29092 18692
rect 28184 18652 29092 18680
rect 27709 18643 27767 18649
rect 29086 18640 29092 18652
rect 29144 18680 29150 18692
rect 29748 18689 29776 18720
rect 29825 18717 29837 18751
rect 29871 18717 29883 18751
rect 30834 18748 30840 18760
rect 30795 18720 30840 18748
rect 29825 18711 29883 18717
rect 30834 18708 30840 18720
rect 30892 18708 30898 18760
rect 31021 18751 31079 18757
rect 31021 18717 31033 18751
rect 31067 18717 31079 18751
rect 31846 18748 31852 18760
rect 31807 18720 31852 18748
rect 31021 18711 31079 18717
rect 29549 18683 29607 18689
rect 29549 18680 29561 18683
rect 29144 18652 29561 18680
rect 29144 18640 29150 18652
rect 29549 18649 29561 18652
rect 29595 18649 29607 18683
rect 29549 18643 29607 18649
rect 29733 18683 29791 18689
rect 29733 18649 29745 18683
rect 29779 18680 29791 18683
rect 30098 18680 30104 18692
rect 29779 18652 30104 18680
rect 29779 18649 29791 18652
rect 29733 18643 29791 18649
rect 30098 18640 30104 18652
rect 30156 18640 30162 18692
rect 31036 18680 31064 18711
rect 31846 18708 31852 18720
rect 31904 18708 31910 18760
rect 32876 18757 32904 18788
rect 33134 18776 33140 18788
rect 33192 18776 33198 18828
rect 35161 18819 35219 18825
rect 35161 18785 35173 18819
rect 35207 18816 35219 18819
rect 35342 18816 35348 18828
rect 35207 18788 35348 18816
rect 35207 18785 35219 18788
rect 35161 18779 35219 18785
rect 35342 18776 35348 18788
rect 35400 18776 35406 18828
rect 32861 18751 32919 18757
rect 32861 18717 32873 18751
rect 32907 18717 32919 18751
rect 32861 18711 32919 18717
rect 33045 18751 33103 18757
rect 33045 18717 33057 18751
rect 33091 18717 33103 18751
rect 33045 18711 33103 18717
rect 32306 18680 32312 18692
rect 31036 18652 32312 18680
rect 32306 18640 32312 18652
rect 32364 18680 32370 18692
rect 33060 18680 33088 18711
rect 33778 18708 33784 18760
rect 33836 18748 33842 18760
rect 35069 18751 35127 18757
rect 35069 18748 35081 18751
rect 33836 18720 35081 18748
rect 33836 18708 33842 18720
rect 35069 18717 35081 18720
rect 35115 18717 35127 18751
rect 36262 18748 36268 18760
rect 36223 18720 36268 18748
rect 35069 18711 35127 18717
rect 36262 18708 36268 18720
rect 36320 18708 36326 18760
rect 36446 18680 36452 18692
rect 32364 18652 33088 18680
rect 36407 18652 36452 18680
rect 32364 18640 32370 18652
rect 36446 18640 36452 18652
rect 36504 18640 36510 18692
rect 38102 18680 38108 18692
rect 38063 18652 38108 18680
rect 38102 18640 38108 18652
rect 38160 18640 38166 18692
rect 23201 18615 23259 18621
rect 23201 18612 23213 18615
rect 22572 18584 23213 18612
rect 17497 18575 17555 18581
rect 23201 18581 23213 18584
rect 23247 18612 23259 18615
rect 23290 18612 23296 18624
rect 23247 18584 23296 18612
rect 23247 18581 23259 18584
rect 23201 18575 23259 18581
rect 23290 18572 23296 18584
rect 23348 18572 23354 18624
rect 26418 18612 26424 18624
rect 26379 18584 26424 18612
rect 26418 18572 26424 18584
rect 26476 18572 26482 18624
rect 26786 18572 26792 18624
rect 26844 18612 26850 18624
rect 27154 18612 27160 18624
rect 26844 18584 27160 18612
rect 26844 18572 26850 18584
rect 27154 18572 27160 18584
rect 27212 18612 27218 18624
rect 27909 18615 27967 18621
rect 27909 18612 27921 18615
rect 27212 18584 27921 18612
rect 27212 18572 27218 18584
rect 27909 18581 27921 18584
rect 27955 18581 27967 18615
rect 28534 18612 28540 18624
rect 28495 18584 28540 18612
rect 27909 18575 27967 18581
rect 28534 18572 28540 18584
rect 28592 18572 28598 18624
rect 30929 18615 30987 18621
rect 30929 18581 30941 18615
rect 30975 18612 30987 18615
rect 31294 18612 31300 18624
rect 30975 18584 31300 18612
rect 30975 18581 30987 18584
rect 30929 18575 30987 18581
rect 31294 18572 31300 18584
rect 31352 18572 31358 18624
rect 31481 18615 31539 18621
rect 31481 18581 31493 18615
rect 31527 18612 31539 18615
rect 31570 18612 31576 18624
rect 31527 18584 31576 18612
rect 31527 18581 31539 18584
rect 31481 18575 31539 18581
rect 31570 18572 31576 18584
rect 31628 18572 31634 18624
rect 32950 18612 32956 18624
rect 32911 18584 32956 18612
rect 32950 18572 32956 18584
rect 33008 18572 33014 18624
rect 34698 18612 34704 18624
rect 34659 18584 34704 18612
rect 34698 18572 34704 18584
rect 34756 18572 34762 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 18138 18368 18144 18420
rect 18196 18408 18202 18420
rect 18417 18411 18475 18417
rect 18417 18408 18429 18411
rect 18196 18380 18429 18408
rect 18196 18368 18202 18380
rect 18417 18377 18429 18380
rect 18463 18377 18475 18411
rect 19334 18408 19340 18420
rect 19295 18380 19340 18408
rect 18417 18371 18475 18377
rect 19334 18368 19340 18380
rect 19392 18368 19398 18420
rect 29825 18411 29883 18417
rect 29825 18377 29837 18411
rect 29871 18408 29883 18411
rect 30098 18408 30104 18420
rect 29871 18380 30104 18408
rect 29871 18377 29883 18380
rect 29825 18371 29883 18377
rect 30098 18368 30104 18380
rect 30156 18368 30162 18420
rect 31481 18411 31539 18417
rect 31481 18377 31493 18411
rect 31527 18408 31539 18411
rect 32214 18408 32220 18420
rect 31527 18380 32220 18408
rect 31527 18377 31539 18380
rect 31481 18371 31539 18377
rect 32214 18368 32220 18380
rect 32272 18408 32278 18420
rect 33134 18408 33140 18420
rect 32272 18380 33140 18408
rect 32272 18368 32278 18380
rect 33134 18368 33140 18380
rect 33192 18368 33198 18420
rect 34238 18368 34244 18420
rect 34296 18408 34302 18420
rect 34333 18411 34391 18417
rect 34333 18408 34345 18411
rect 34296 18380 34345 18408
rect 34296 18368 34302 18380
rect 34333 18377 34345 18380
rect 34379 18377 34391 18411
rect 34333 18371 34391 18377
rect 36446 18368 36452 18420
rect 36504 18408 36510 18420
rect 37553 18411 37611 18417
rect 37553 18408 37565 18411
rect 36504 18380 37565 18408
rect 36504 18368 36510 18380
rect 37553 18377 37565 18380
rect 37599 18377 37611 18411
rect 37553 18371 37611 18377
rect 7374 18300 7380 18352
rect 7432 18340 7438 18352
rect 8110 18340 8116 18352
rect 7432 18312 8116 18340
rect 7432 18300 7438 18312
rect 8110 18300 8116 18312
rect 8168 18340 8174 18352
rect 8168 18312 37504 18340
rect 8168 18300 8174 18312
rect 37476 18284 37504 18312
rect 17034 18272 17040 18284
rect 16995 18244 17040 18272
rect 17034 18232 17040 18244
rect 17092 18232 17098 18284
rect 17310 18281 17316 18284
rect 17304 18272 17316 18281
rect 17271 18244 17316 18272
rect 17304 18235 17316 18244
rect 17310 18232 17316 18235
rect 17368 18232 17374 18284
rect 19426 18232 19432 18284
rect 19484 18272 19490 18284
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 19484 18244 19625 18272
rect 19484 18232 19490 18244
rect 19613 18241 19625 18244
rect 19659 18241 19671 18275
rect 28442 18272 28448 18284
rect 28403 18244 28448 18272
rect 19613 18235 19671 18241
rect 28442 18232 28448 18244
rect 28500 18232 28506 18284
rect 28534 18232 28540 18284
rect 28592 18272 28598 18284
rect 28701 18275 28759 18281
rect 28701 18272 28713 18275
rect 28592 18244 28713 18272
rect 28592 18232 28598 18244
rect 28701 18241 28713 18244
rect 28747 18241 28759 18275
rect 31294 18272 31300 18284
rect 31255 18244 31300 18272
rect 28701 18235 28759 18241
rect 31294 18232 31300 18244
rect 31352 18232 31358 18284
rect 31570 18232 31576 18284
rect 31628 18272 31634 18284
rect 31628 18244 31673 18272
rect 31628 18232 31634 18244
rect 32674 18232 32680 18284
rect 32732 18272 32738 18284
rect 33226 18281 33232 18284
rect 32953 18275 33011 18281
rect 32953 18272 32965 18275
rect 32732 18244 32965 18272
rect 32732 18232 32738 18244
rect 32953 18241 32965 18244
rect 32999 18241 33011 18275
rect 32953 18235 33011 18241
rect 33220 18235 33232 18281
rect 33284 18272 33290 18284
rect 33284 18244 33320 18272
rect 33226 18232 33232 18235
rect 33284 18232 33290 18244
rect 36262 18232 36268 18284
rect 36320 18272 36326 18284
rect 36541 18275 36599 18281
rect 36541 18272 36553 18275
rect 36320 18244 36553 18272
rect 36320 18232 36326 18244
rect 36541 18241 36553 18244
rect 36587 18241 36599 18275
rect 37458 18272 37464 18284
rect 37371 18244 37464 18272
rect 36541 18235 36599 18241
rect 37458 18232 37464 18244
rect 37516 18232 37522 18284
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18173 19395 18207
rect 19337 18167 19395 18173
rect 19521 18207 19579 18213
rect 19521 18173 19533 18207
rect 19567 18204 19579 18207
rect 19978 18204 19984 18216
rect 19567 18176 19984 18204
rect 19567 18173 19579 18176
rect 19521 18167 19579 18173
rect 19352 18136 19380 18167
rect 19978 18164 19984 18176
rect 20036 18164 20042 18216
rect 31110 18164 31116 18216
rect 31168 18204 31174 18216
rect 31205 18207 31263 18213
rect 31205 18204 31217 18207
rect 31168 18176 31217 18204
rect 31168 18164 31174 18176
rect 31205 18173 31217 18176
rect 31251 18204 31263 18207
rect 32766 18204 32772 18216
rect 31251 18176 32772 18204
rect 31251 18173 31263 18176
rect 31205 18167 31263 18173
rect 32766 18164 32772 18176
rect 32824 18164 32830 18216
rect 20162 18136 20168 18148
rect 19352 18108 20168 18136
rect 20162 18096 20168 18108
rect 20220 18096 20226 18148
rect 1670 18068 1676 18080
rect 1631 18040 1676 18068
rect 1670 18028 1676 18040
rect 1728 18028 1734 18080
rect 31202 18068 31208 18080
rect 31163 18040 31208 18068
rect 31202 18028 31208 18040
rect 31260 18028 31266 18080
rect 36078 18068 36084 18080
rect 36039 18040 36084 18068
rect 36078 18028 36084 18040
rect 36136 18028 36142 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 27157 17867 27215 17873
rect 27157 17833 27169 17867
rect 27203 17864 27215 17867
rect 27246 17864 27252 17876
rect 27203 17836 27252 17864
rect 27203 17833 27215 17836
rect 27157 17827 27215 17833
rect 27246 17824 27252 17836
rect 27304 17824 27310 17876
rect 30193 17867 30251 17873
rect 30193 17833 30205 17867
rect 30239 17864 30251 17867
rect 30834 17864 30840 17876
rect 30239 17836 30840 17864
rect 30239 17833 30251 17836
rect 30193 17827 30251 17833
rect 30834 17824 30840 17836
rect 30892 17824 30898 17876
rect 32950 17824 32956 17876
rect 33008 17864 33014 17876
rect 33045 17867 33103 17873
rect 33045 17864 33057 17867
rect 33008 17836 33057 17864
rect 33008 17824 33014 17836
rect 33045 17833 33057 17836
rect 33091 17833 33103 17867
rect 33045 17827 33103 17833
rect 32861 17799 32919 17805
rect 32861 17765 32873 17799
rect 32907 17796 32919 17799
rect 33226 17796 33232 17808
rect 32907 17768 33232 17796
rect 32907 17765 32919 17768
rect 32861 17759 32919 17765
rect 33226 17756 33232 17768
rect 33284 17756 33290 17808
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 1670 17728 1676 17740
rect 1443 17700 1676 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 1670 17688 1676 17700
rect 1728 17688 1734 17740
rect 2774 17728 2780 17740
rect 2735 17700 2780 17728
rect 2774 17688 2780 17700
rect 2832 17688 2838 17740
rect 25038 17688 25044 17740
rect 25096 17728 25102 17740
rect 25777 17731 25835 17737
rect 25777 17728 25789 17731
rect 25096 17700 25789 17728
rect 25096 17688 25102 17700
rect 25777 17697 25789 17700
rect 25823 17697 25835 17731
rect 25777 17691 25835 17697
rect 31573 17731 31631 17737
rect 31573 17697 31585 17731
rect 31619 17728 31631 17731
rect 32674 17728 32680 17740
rect 31619 17700 32680 17728
rect 31619 17697 31631 17700
rect 31573 17691 31631 17697
rect 32674 17688 32680 17700
rect 32732 17688 32738 17740
rect 32766 17688 32772 17740
rect 32824 17728 32830 17740
rect 32953 17731 33011 17737
rect 32953 17728 32965 17731
rect 32824 17700 32965 17728
rect 32824 17688 32830 17700
rect 32953 17697 32965 17700
rect 32999 17697 33011 17731
rect 32953 17691 33011 17697
rect 36078 17688 36084 17740
rect 36136 17728 36142 17740
rect 36265 17731 36323 17737
rect 36265 17728 36277 17731
rect 36136 17700 36277 17728
rect 36136 17688 36142 17700
rect 36265 17697 36277 17700
rect 36311 17697 36323 17731
rect 38102 17728 38108 17740
rect 38063 17700 38108 17728
rect 36265 17691 36323 17697
rect 38102 17688 38108 17700
rect 38160 17688 38166 17740
rect 26044 17663 26102 17669
rect 26044 17629 26056 17663
rect 26090 17660 26102 17663
rect 26418 17660 26424 17672
rect 26090 17632 26424 17660
rect 26090 17629 26102 17632
rect 26044 17623 26102 17629
rect 26418 17620 26424 17632
rect 26476 17620 26482 17672
rect 33134 17660 33140 17672
rect 33095 17632 33140 17660
rect 33134 17620 33140 17632
rect 33192 17620 33198 17672
rect 33321 17663 33379 17669
rect 33321 17629 33333 17663
rect 33367 17660 33379 17663
rect 34698 17660 34704 17672
rect 33367 17632 34704 17660
rect 33367 17629 33379 17632
rect 33321 17623 33379 17629
rect 34698 17620 34704 17632
rect 34756 17620 34762 17672
rect 1581 17595 1639 17601
rect 1581 17561 1593 17595
rect 1627 17592 1639 17595
rect 2130 17592 2136 17604
rect 1627 17564 2136 17592
rect 1627 17561 1639 17564
rect 1581 17555 1639 17561
rect 2130 17552 2136 17564
rect 2188 17552 2194 17604
rect 31202 17552 31208 17604
rect 31260 17592 31266 17604
rect 31306 17595 31364 17601
rect 31306 17592 31318 17595
rect 31260 17564 31318 17592
rect 31260 17552 31266 17564
rect 31306 17561 31318 17564
rect 31352 17561 31364 17595
rect 36446 17592 36452 17604
rect 36407 17564 36452 17592
rect 31306 17555 31364 17561
rect 36446 17552 36452 17564
rect 36504 17552 36510 17604
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 2130 17320 2136 17332
rect 2091 17292 2136 17320
rect 2130 17280 2136 17292
rect 2188 17280 2194 17332
rect 36446 17280 36452 17332
rect 36504 17320 36510 17332
rect 37553 17323 37611 17329
rect 37553 17320 37565 17323
rect 36504 17292 37565 17320
rect 36504 17280 36510 17292
rect 37553 17289 37565 17292
rect 37599 17289 37611 17323
rect 37553 17283 37611 17289
rect 2222 17184 2228 17196
rect 2135 17156 2228 17184
rect 2222 17144 2228 17156
rect 2280 17184 2286 17196
rect 15378 17184 15384 17196
rect 2280 17156 15384 17184
rect 2280 17144 2286 17156
rect 15378 17144 15384 17156
rect 15436 17184 15442 17196
rect 15562 17184 15568 17196
rect 15436 17156 15568 17184
rect 15436 17144 15442 17156
rect 15562 17144 15568 17156
rect 15620 17144 15626 17196
rect 37458 17184 37464 17196
rect 37419 17156 37464 17184
rect 37458 17144 37464 17156
rect 37516 17184 37522 17196
rect 37642 17184 37648 17196
rect 37516 17156 37648 17184
rect 37516 17144 37522 17156
rect 37642 17144 37648 17156
rect 37700 17144 37706 17196
rect 1394 16980 1400 16992
rect 1355 16952 1400 16980
rect 1394 16940 1400 16952
rect 1452 16940 1458 16992
rect 36262 16940 36268 16992
rect 36320 16980 36326 16992
rect 36541 16983 36599 16989
rect 36541 16980 36553 16983
rect 36320 16952 36553 16980
rect 36320 16940 36326 16952
rect 36541 16949 36553 16952
rect 36587 16949 36599 16983
rect 36541 16943 36599 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 1394 16640 1400 16652
rect 1355 16612 1400 16640
rect 1394 16600 1400 16612
rect 1452 16600 1458 16652
rect 1854 16640 1860 16652
rect 1815 16612 1860 16640
rect 1854 16600 1860 16612
rect 1912 16600 1918 16652
rect 36262 16640 36268 16652
rect 36223 16612 36268 16640
rect 36262 16600 36268 16612
rect 36320 16600 36326 16652
rect 38102 16640 38108 16652
rect 38063 16612 38108 16640
rect 38102 16600 38108 16612
rect 38160 16600 38166 16652
rect 1581 16507 1639 16513
rect 1581 16473 1593 16507
rect 1627 16504 1639 16507
rect 2038 16504 2044 16516
rect 1627 16476 2044 16504
rect 1627 16473 1639 16476
rect 1581 16467 1639 16473
rect 2038 16464 2044 16476
rect 2096 16464 2102 16516
rect 36446 16504 36452 16516
rect 36407 16476 36452 16504
rect 36446 16464 36452 16476
rect 36504 16464 36510 16516
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 2038 16232 2044 16244
rect 1999 16204 2044 16232
rect 2038 16192 2044 16204
rect 2096 16192 2102 16244
rect 36446 16192 36452 16244
rect 36504 16232 36510 16244
rect 37553 16235 37611 16241
rect 37553 16232 37565 16235
rect 36504 16204 37565 16232
rect 36504 16192 36510 16204
rect 37553 16201 37565 16204
rect 37599 16201 37611 16235
rect 37553 16195 37611 16201
rect 2130 16096 2136 16108
rect 2091 16068 2136 16096
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 37458 16096 37464 16108
rect 37419 16068 37464 16096
rect 37458 16056 37464 16068
rect 37516 16096 37522 16108
rect 38010 16096 38016 16108
rect 37516 16068 38016 16096
rect 37516 16056 37522 16068
rect 38010 16056 38016 16068
rect 38068 16056 38074 16108
rect 2777 15895 2835 15901
rect 2777 15861 2789 15895
rect 2823 15892 2835 15895
rect 3234 15892 3240 15904
rect 2823 15864 3240 15892
rect 2823 15861 2835 15864
rect 2777 15855 2835 15861
rect 3234 15852 3240 15864
rect 3292 15852 3298 15904
rect 36262 15852 36268 15904
rect 36320 15892 36326 15904
rect 36541 15895 36599 15901
rect 36541 15892 36553 15895
rect 36320 15864 36553 15892
rect 36320 15852 36326 15864
rect 36541 15861 36553 15864
rect 36587 15861 36599 15895
rect 36541 15855 36599 15861
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 1394 15552 1400 15564
rect 1355 15524 1400 15552
rect 1394 15512 1400 15524
rect 1452 15512 1458 15564
rect 3234 15552 3240 15564
rect 3195 15524 3240 15552
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 36262 15552 36268 15564
rect 36223 15524 36268 15552
rect 36262 15512 36268 15524
rect 36320 15512 36326 15564
rect 38102 15552 38108 15564
rect 38063 15524 38108 15552
rect 38102 15512 38108 15524
rect 38160 15512 38166 15564
rect 3050 15416 3056 15428
rect 3011 15388 3056 15416
rect 3050 15376 3056 15388
rect 3108 15376 3114 15428
rect 36446 15416 36452 15428
rect 36407 15388 36452 15416
rect 36446 15376 36452 15388
rect 36504 15376 36510 15428
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 1949 15147 2007 15153
rect 1949 15113 1961 15147
rect 1995 15144 2007 15147
rect 3050 15144 3056 15156
rect 1995 15116 3056 15144
rect 1995 15113 2007 15116
rect 1949 15107 2007 15113
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 36446 15104 36452 15156
rect 36504 15144 36510 15156
rect 36541 15147 36599 15153
rect 36541 15144 36553 15147
rect 36504 15116 36553 15144
rect 36504 15104 36510 15116
rect 36541 15113 36553 15116
rect 36587 15113 36599 15147
rect 36541 15107 36599 15113
rect 1857 15011 1915 15017
rect 1857 14977 1869 15011
rect 1903 15008 1915 15011
rect 2314 15008 2320 15020
rect 1903 14980 2320 15008
rect 1903 14977 1915 14980
rect 1857 14971 1915 14977
rect 2314 14968 2320 14980
rect 2372 15008 2378 15020
rect 14458 15008 14464 15020
rect 2372 14980 14464 15008
rect 2372 14968 2378 14980
rect 14458 14968 14464 14980
rect 14516 15008 14522 15020
rect 36354 15008 36360 15020
rect 14516 14980 36360 15008
rect 14516 14968 14522 14980
rect 36354 14968 36360 14980
rect 36412 15008 36418 15020
rect 36449 15011 36507 15017
rect 36449 15008 36461 15011
rect 36412 14980 36461 15008
rect 36412 14968 36418 14980
rect 36449 14977 36461 14980
rect 36495 14977 36507 15011
rect 36449 14971 36507 14977
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1670 14356 1676 14408
rect 1728 14396 1734 14408
rect 1765 14399 1823 14405
rect 1765 14396 1777 14399
rect 1728 14368 1777 14396
rect 1728 14356 1734 14368
rect 1765 14365 1777 14368
rect 1811 14365 1823 14399
rect 1765 14359 1823 14365
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 1854 13852 1860 13864
rect 1815 13824 1860 13852
rect 1854 13812 1860 13824
rect 1912 13812 1918 13864
rect 2774 13852 2780 13864
rect 2735 13824 2780 13852
rect 2774 13812 2780 13824
rect 2832 13812 2838 13864
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 1854 13472 1860 13524
rect 1912 13512 1918 13524
rect 2133 13515 2191 13521
rect 2133 13512 2145 13515
rect 1912 13484 2145 13512
rect 1912 13472 1918 13484
rect 2133 13481 2145 13484
rect 2179 13481 2191 13515
rect 2133 13475 2191 13481
rect 1581 13311 1639 13317
rect 1581 13277 1593 13311
rect 1627 13308 1639 13311
rect 1670 13308 1676 13320
rect 1627 13280 1676 13308
rect 1627 13277 1639 13280
rect 1581 13271 1639 13277
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 2222 13308 2228 13320
rect 2183 13280 2228 13308
rect 2222 13268 2228 13280
rect 2280 13268 2286 13320
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 37826 12900 37832 12912
rect 37787 12872 37832 12900
rect 37826 12860 37832 12872
rect 37884 12860 37890 12912
rect 1670 12832 1676 12844
rect 1631 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 38102 12832 38108 12844
rect 38063 12804 38108 12832
rect 38102 12792 38108 12804
rect 38160 12792 38166 12844
rect 1854 12764 1860 12776
rect 1815 12736 1860 12764
rect 1854 12724 1860 12736
rect 1912 12724 1918 12776
rect 2774 12764 2780 12776
rect 2735 12736 2780 12764
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 1854 12384 1860 12436
rect 1912 12424 1918 12436
rect 2133 12427 2191 12433
rect 2133 12424 2145 12427
rect 1912 12396 2145 12424
rect 1912 12384 1918 12396
rect 2133 12393 2145 12396
rect 2179 12393 2191 12427
rect 2133 12387 2191 12393
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 9398 12220 9404 12232
rect 2271 12192 9404 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 37829 12223 37887 12229
rect 37829 12189 37841 12223
rect 37875 12220 37887 12223
rect 38102 12220 38108 12232
rect 37875 12192 38108 12220
rect 37875 12189 37887 12192
rect 37829 12183 37887 12189
rect 38102 12180 38108 12192
rect 38160 12180 38166 12232
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 8754 11704 8760 11756
rect 8812 11744 8818 11756
rect 37366 11744 37372 11756
rect 8812 11716 37372 11744
rect 8812 11704 8818 11716
rect 37366 11704 37372 11716
rect 37424 11704 37430 11756
rect 37461 11543 37519 11549
rect 37461 11509 37473 11543
rect 37507 11540 37519 11543
rect 37918 11540 37924 11552
rect 37507 11512 37924 11540
rect 37507 11509 37519 11512
rect 37461 11503 37519 11509
rect 37918 11500 37924 11512
rect 37976 11500 37982 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 37182 11200 37188 11212
rect 37143 11172 37188 11200
rect 37182 11160 37188 11172
rect 37240 11160 37246 11212
rect 37918 11200 37924 11212
rect 37879 11172 37924 11200
rect 37918 11160 37924 11172
rect 37976 11160 37982 11212
rect 38102 11200 38108 11212
rect 38063 11172 38108 11200
rect 38102 11160 38108 11172
rect 38160 11160 38166 11212
rect 2041 11135 2099 11141
rect 2041 11101 2053 11135
rect 2087 11132 2099 11135
rect 2130 11132 2136 11144
rect 2087 11104 2136 11132
rect 2087 11101 2099 11104
rect 2041 11095 2099 11101
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 3418 11132 3424 11144
rect 2731 11104 3424 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 1949 11067 2007 11073
rect 1949 11033 1961 11067
rect 1995 11064 2007 11067
rect 3234 11064 3240 11076
rect 1995 11036 3240 11064
rect 1995 11033 2007 11036
rect 1949 11027 2007 11033
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 3234 10724 3240 10736
rect 3195 10696 3240 10724
rect 3234 10684 3240 10696
rect 3292 10684 3298 10736
rect 3418 10616 3424 10668
rect 3476 10656 3482 10668
rect 37461 10659 37519 10665
rect 3476 10628 3521 10656
rect 3476 10616 3482 10628
rect 37461 10625 37473 10659
rect 37507 10656 37519 10659
rect 37550 10656 37556 10668
rect 37507 10628 37556 10656
rect 37507 10625 37519 10628
rect 37461 10619 37519 10625
rect 37550 10616 37556 10628
rect 37608 10616 37614 10668
rect 1578 10588 1584 10600
rect 1539 10560 1584 10588
rect 1578 10548 1584 10560
rect 1636 10548 1642 10600
rect 36446 10412 36452 10464
rect 36504 10452 36510 10464
rect 37369 10455 37427 10461
rect 37369 10452 37381 10455
rect 36504 10424 37381 10452
rect 36504 10412 36510 10424
rect 37369 10421 37381 10424
rect 37415 10421 37427 10455
rect 38102 10452 38108 10464
rect 38063 10424 38108 10452
rect 37369 10415 37427 10421
rect 38102 10412 38108 10424
rect 38160 10412 38166 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 36446 10112 36452 10124
rect 36407 10084 36452 10112
rect 36446 10072 36452 10084
rect 36504 10072 36510 10124
rect 1854 10044 1860 10056
rect 1815 10016 1860 10044
rect 1854 10004 1860 10016
rect 1912 10004 1918 10056
rect 2498 10044 2504 10056
rect 2459 10016 2504 10044
rect 2498 10004 2504 10016
rect 2556 10044 2562 10056
rect 20346 10044 20352 10056
rect 2556 10016 20352 10044
rect 2556 10004 2562 10016
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 36262 10044 36268 10056
rect 36223 10016 36268 10044
rect 36262 10004 36268 10016
rect 36320 10004 36326 10056
rect 38010 9936 38016 9988
rect 38068 9976 38074 9988
rect 38105 9979 38163 9985
rect 38105 9976 38117 9979
rect 38068 9948 38117 9976
rect 38068 9936 38074 9948
rect 38105 9945 38117 9948
rect 38151 9945 38163 9979
rect 38105 9939 38163 9945
rect 2038 9868 2044 9920
rect 2096 9908 2102 9920
rect 2409 9911 2467 9917
rect 2409 9908 2421 9911
rect 2096 9880 2421 9908
rect 2096 9868 2102 9880
rect 2409 9877 2421 9880
rect 2455 9877 2467 9911
rect 2409 9871 2467 9877
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 2038 9636 2044 9648
rect 1999 9608 2044 9636
rect 2038 9596 2044 9608
rect 2096 9596 2102 9648
rect 1854 9568 1860 9580
rect 1815 9540 1860 9568
rect 1854 9528 1860 9540
rect 1912 9528 1918 9580
rect 36262 9528 36268 9580
rect 36320 9568 36326 9580
rect 36541 9571 36599 9577
rect 36541 9568 36553 9571
rect 36320 9540 36553 9568
rect 36320 9528 36326 9540
rect 36541 9537 36553 9540
rect 36587 9537 36599 9571
rect 37458 9568 37464 9580
rect 37419 9540 37464 9568
rect 36541 9531 36599 9537
rect 37458 9528 37464 9540
rect 37516 9528 37522 9580
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 2832 9472 2877 9500
rect 2832 9460 2838 9472
rect 37553 9367 37611 9373
rect 37553 9333 37565 9367
rect 37599 9364 37611 9367
rect 37918 9364 37924 9376
rect 37599 9336 37924 9364
rect 37599 9333 37611 9336
rect 37553 9327 37611 9333
rect 37918 9324 37924 9336
rect 37976 9324 37982 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 37182 9024 37188 9036
rect 37143 8996 37188 9024
rect 37182 8984 37188 8996
rect 37240 8984 37246 9036
rect 37918 9024 37924 9036
rect 37879 8996 37924 9024
rect 37918 8984 37924 8996
rect 37976 8984 37982 9036
rect 38102 9024 38108 9036
rect 38063 8996 38108 9024
rect 38102 8984 38108 8996
rect 38160 8984 38166 9036
rect 2038 8956 2044 8968
rect 1999 8928 2044 8956
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 2866 8956 2872 8968
rect 2731 8928 2872 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 2593 8823 2651 8829
rect 2593 8820 2605 8823
rect 2280 8792 2605 8820
rect 2280 8780 2286 8792
rect 2593 8789 2605 8792
rect 2639 8789 2651 8823
rect 2593 8783 2651 8789
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 2222 8548 2228 8560
rect 2183 8520 2228 8548
rect 2222 8508 2228 8520
rect 2280 8508 2286 8560
rect 2038 8480 2044 8492
rect 1999 8452 2044 8480
rect 2038 8440 2044 8452
rect 2096 8440 2102 8492
rect 2866 8412 2872 8424
rect 2827 8384 2872 8412
rect 2866 8372 2872 8384
rect 2924 8372 2930 8424
rect 37829 8347 37887 8353
rect 37829 8313 37841 8347
rect 37875 8344 37887 8347
rect 38102 8344 38108 8356
rect 37875 8316 38108 8344
rect 37875 8313 37887 8316
rect 37829 8307 37887 8313
rect 38102 8304 38108 8316
rect 38160 8304 38166 8356
rect 1394 8276 1400 8288
rect 1355 8248 1400 8276
rect 1394 8236 1400 8248
rect 1452 8236 1458 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1394 7936 1400 7948
rect 1355 7908 1400 7936
rect 1394 7896 1400 7908
rect 1452 7896 1458 7948
rect 2774 7896 2780 7948
rect 2832 7936 2838 7948
rect 2832 7908 2877 7936
rect 2832 7896 2838 7908
rect 37826 7868 37832 7880
rect 37787 7840 37832 7868
rect 37826 7828 37832 7840
rect 37884 7828 37890 7880
rect 1581 7803 1639 7809
rect 1581 7769 1593 7803
rect 1627 7800 1639 7803
rect 2222 7800 2228 7812
rect 1627 7772 2228 7800
rect 1627 7769 1639 7772
rect 1581 7763 1639 7769
rect 2222 7760 2228 7772
rect 2280 7760 2286 7812
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 2222 7528 2228 7540
rect 2183 7500 2228 7528
rect 2222 7488 2228 7500
rect 2280 7488 2286 7540
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 7006 7392 7012 7404
rect 2363 7364 7012 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 7006 7352 7012 7364
rect 7064 7352 7070 7404
rect 37461 7395 37519 7401
rect 37461 7361 37473 7395
rect 37507 7392 37519 7395
rect 37642 7392 37648 7404
rect 37507 7364 37648 7392
rect 37507 7361 37519 7364
rect 37461 7355 37519 7361
rect 37642 7352 37648 7364
rect 37700 7352 37706 7404
rect 1394 7148 1400 7200
rect 1452 7188 1458 7200
rect 1489 7191 1547 7197
rect 1489 7188 1501 7191
rect 1452 7160 1501 7188
rect 1452 7148 1458 7160
rect 1489 7157 1501 7160
rect 1535 7157 1547 7191
rect 1489 7151 1547 7157
rect 37553 7191 37611 7197
rect 37553 7157 37565 7191
rect 37599 7188 37611 7191
rect 37918 7188 37924 7200
rect 37599 7160 37924 7188
rect 37599 7157 37611 7160
rect 37553 7151 37611 7157
rect 37918 7148 37924 7160
rect 37976 7148 37982 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1394 6848 1400 6860
rect 1355 6820 1400 6848
rect 1394 6808 1400 6820
rect 1452 6808 1458 6860
rect 2774 6808 2780 6860
rect 2832 6848 2838 6860
rect 37182 6848 37188 6860
rect 2832 6820 2877 6848
rect 37143 6820 37188 6848
rect 2832 6808 2838 6820
rect 37182 6808 37188 6820
rect 37240 6808 37246 6860
rect 37918 6848 37924 6860
rect 37879 6820 37924 6848
rect 37918 6808 37924 6820
rect 37976 6808 37982 6860
rect 38102 6848 38108 6860
rect 38063 6820 38108 6848
rect 38102 6808 38108 6820
rect 38160 6808 38166 6860
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 2038 6712 2044 6724
rect 1627 6684 2044 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 2038 6672 2044 6684
rect 2096 6672 2102 6724
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 2038 6440 2044 6452
rect 1999 6412 2044 6440
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 2130 6304 2136 6316
rect 2091 6276 2136 6304
rect 2130 6264 2136 6276
rect 2188 6304 2194 6316
rect 2406 6304 2412 6316
rect 2188 6276 2412 6304
rect 2188 6264 2194 6276
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 37461 6307 37519 6313
rect 37461 6273 37473 6307
rect 37507 6304 37519 6307
rect 37550 6304 37556 6316
rect 37507 6276 37556 6304
rect 37507 6273 37519 6276
rect 37461 6267 37519 6273
rect 37550 6264 37556 6276
rect 37608 6264 37614 6316
rect 35342 6236 35348 6248
rect 35303 6208 35348 6236
rect 35342 6196 35348 6208
rect 35400 6196 35406 6248
rect 36538 6236 36544 6248
rect 36499 6208 36544 6236
rect 36538 6196 36544 6208
rect 36596 6196 36602 6248
rect 36725 6239 36783 6245
rect 36725 6205 36737 6239
rect 36771 6236 36783 6239
rect 37826 6236 37832 6248
rect 36771 6208 37832 6236
rect 36771 6205 36783 6208
rect 36725 6199 36783 6205
rect 37826 6196 37832 6208
rect 37884 6196 37890 6248
rect 2777 6103 2835 6109
rect 2777 6069 2789 6103
rect 2823 6100 2835 6103
rect 3234 6100 3240 6112
rect 2823 6072 3240 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 3234 6060 3240 6072
rect 3292 6060 3298 6112
rect 37553 6103 37611 6109
rect 37553 6069 37565 6103
rect 37599 6100 37611 6103
rect 37918 6100 37924 6112
rect 37599 6072 37924 6100
rect 37599 6069 37611 6072
rect 37553 6063 37611 6069
rect 37918 6060 37924 6072
rect 37976 6060 37982 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 37734 5788 37740 5840
rect 37792 5828 37798 5840
rect 37792 5800 38148 5828
rect 37792 5788 37798 5800
rect 3234 5760 3240 5772
rect 3195 5732 3240 5760
rect 3234 5720 3240 5732
rect 3292 5720 3298 5772
rect 37182 5760 37188 5772
rect 37143 5732 37188 5760
rect 37182 5720 37188 5732
rect 37240 5720 37246 5772
rect 37918 5760 37924 5772
rect 37879 5732 37924 5760
rect 37918 5720 37924 5732
rect 37976 5720 37982 5772
rect 38120 5769 38148 5800
rect 38105 5763 38163 5769
rect 38105 5729 38117 5763
rect 38151 5729 38163 5763
rect 38105 5723 38163 5729
rect 33410 5692 33416 5704
rect 33371 5664 33416 5692
rect 33410 5652 33416 5664
rect 33468 5652 33474 5704
rect 34514 5652 34520 5704
rect 34572 5692 34578 5704
rect 34885 5695 34943 5701
rect 34885 5692 34897 5695
rect 34572 5664 34897 5692
rect 34572 5652 34578 5664
rect 34885 5661 34897 5664
rect 34931 5661 34943 5695
rect 34885 5655 34943 5661
rect 35713 5695 35771 5701
rect 35713 5661 35725 5695
rect 35759 5692 35771 5695
rect 36446 5692 36452 5704
rect 35759 5664 36452 5692
rect 35759 5661 35771 5664
rect 35713 5655 35771 5661
rect 36446 5652 36452 5664
rect 36504 5652 36510 5704
rect 1394 5624 1400 5636
rect 1355 5596 1400 5624
rect 1394 5584 1400 5596
rect 1452 5584 1458 5636
rect 3050 5624 3056 5636
rect 3011 5596 3056 5624
rect 3050 5584 3056 5596
rect 3108 5584 3114 5636
rect 35526 5516 35532 5568
rect 35584 5556 35590 5568
rect 35621 5559 35679 5565
rect 35621 5556 35633 5559
rect 35584 5528 35633 5556
rect 35584 5516 35590 5528
rect 35621 5525 35633 5528
rect 35667 5525 35679 5559
rect 35621 5519 35679 5525
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 3050 5352 3056 5364
rect 1995 5324 3056 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 36265 5355 36323 5361
rect 36265 5321 36277 5355
rect 36311 5352 36323 5355
rect 36538 5352 36544 5364
rect 36311 5324 36544 5352
rect 36311 5321 36323 5324
rect 36265 5315 36323 5321
rect 36538 5312 36544 5324
rect 36596 5312 36602 5364
rect 14550 5244 14556 5296
rect 14608 5284 14614 5296
rect 35250 5284 35256 5296
rect 14608 5256 34836 5284
rect 35211 5256 35256 5284
rect 14608 5244 14614 5256
rect 2041 5219 2099 5225
rect 2041 5185 2053 5219
rect 2087 5216 2099 5219
rect 2314 5216 2320 5228
rect 2087 5188 2320 5216
rect 2087 5185 2099 5188
rect 2041 5179 2099 5185
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 32674 5216 32680 5228
rect 32635 5188 32680 5216
rect 32674 5176 32680 5188
rect 32732 5176 32738 5228
rect 33410 5216 33416 5228
rect 33371 5188 33416 5216
rect 33410 5176 33416 5188
rect 33468 5176 33474 5228
rect 34808 5216 34836 5256
rect 35250 5244 35256 5256
rect 35308 5244 35314 5296
rect 36357 5219 36415 5225
rect 36357 5216 36369 5219
rect 34808 5188 36369 5216
rect 36357 5185 36369 5188
rect 36403 5216 36415 5219
rect 37277 5219 37335 5225
rect 37277 5216 37289 5219
rect 36403 5188 37289 5216
rect 36403 5185 36415 5188
rect 36357 5179 36415 5185
rect 37277 5185 37289 5188
rect 37323 5185 37335 5219
rect 37277 5179 37335 5185
rect 37826 5176 37832 5228
rect 37884 5216 37890 5228
rect 37921 5219 37979 5225
rect 37921 5216 37933 5219
rect 37884 5188 37933 5216
rect 37884 5176 37890 5188
rect 37921 5185 37933 5188
rect 37967 5185 37979 5219
rect 37921 5179 37979 5185
rect 2958 5148 2964 5160
rect 2919 5120 2964 5148
rect 2958 5108 2964 5120
rect 3016 5108 3022 5160
rect 3145 5151 3203 5157
rect 3145 5117 3157 5151
rect 3191 5148 3203 5151
rect 3878 5148 3884 5160
rect 3191 5120 3884 5148
rect 3191 5117 3203 5120
rect 3145 5111 3203 5117
rect 3878 5108 3884 5120
rect 3936 5108 3942 5160
rect 3970 5108 3976 5160
rect 4028 5148 4034 5160
rect 32769 5151 32827 5157
rect 4028 5120 4073 5148
rect 4028 5108 4034 5120
rect 32769 5117 32781 5151
rect 32815 5148 32827 5151
rect 33597 5151 33655 5157
rect 33597 5148 33609 5151
rect 32815 5120 33609 5148
rect 32815 5117 32827 5120
rect 32769 5111 32827 5117
rect 33597 5117 33609 5120
rect 33643 5117 33655 5151
rect 33597 5111 33655 5117
rect 33962 5040 33968 5092
rect 34020 5080 34026 5092
rect 37369 5083 37427 5089
rect 37369 5080 37381 5083
rect 34020 5052 37381 5080
rect 34020 5040 34026 5052
rect 37369 5049 37381 5052
rect 37415 5049 37427 5083
rect 37369 5043 37427 5049
rect 6362 5012 6368 5024
rect 6323 4984 6368 5012
rect 6362 4972 6368 4984
rect 6420 4972 6426 5024
rect 7469 5015 7527 5021
rect 7469 4981 7481 5015
rect 7515 5012 7527 5015
rect 8938 5012 8944 5024
rect 7515 4984 8944 5012
rect 7515 4981 7527 4984
rect 7469 4975 7527 4981
rect 8938 4972 8944 4984
rect 8996 4972 9002 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 2958 4808 2964 4820
rect 2919 4780 2964 4808
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 3878 4808 3884 4820
rect 3839 4780 3884 4808
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 4062 4700 4068 4752
rect 4120 4740 4126 4752
rect 34606 4740 34612 4752
rect 4120 4712 6868 4740
rect 4120 4700 4126 4712
rect 5261 4675 5319 4681
rect 5261 4641 5273 4675
rect 5307 4672 5319 4675
rect 6178 4672 6184 4684
rect 5307 4644 6184 4672
rect 5307 4641 5319 4644
rect 5261 4635 5319 4641
rect 6178 4632 6184 4644
rect 6236 4632 6242 4684
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 6840 4681 6868 4712
rect 33704 4712 34612 4740
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4641 6883 4675
rect 6825 4635 6883 4641
rect 15470 4632 15476 4684
rect 15528 4672 15534 4684
rect 33704 4681 33732 4712
rect 34606 4700 34612 4712
rect 34664 4700 34670 4752
rect 15657 4675 15715 4681
rect 15657 4672 15669 4675
rect 15528 4644 15669 4672
rect 15528 4632 15534 4644
rect 15657 4641 15669 4644
rect 15703 4641 15715 4675
rect 15657 4635 15715 4641
rect 33689 4675 33747 4681
rect 33689 4641 33701 4675
rect 33735 4641 33747 4675
rect 33962 4672 33968 4684
rect 33923 4644 33968 4672
rect 33689 4635 33747 4641
rect 33962 4632 33968 4644
rect 34020 4632 34026 4684
rect 34149 4675 34207 4681
rect 34149 4641 34161 4675
rect 34195 4672 34207 4675
rect 34514 4672 34520 4684
rect 34195 4644 34520 4672
rect 34195 4641 34207 4644
rect 34149 4635 34207 4641
rect 34514 4632 34520 4644
rect 34572 4632 34578 4684
rect 35526 4672 35532 4684
rect 35487 4644 35532 4672
rect 35526 4632 35532 4644
rect 35584 4632 35590 4684
rect 36078 4672 36084 4684
rect 36039 4644 36084 4672
rect 36078 4632 36084 4644
rect 36136 4632 36142 4684
rect 1394 4564 1400 4616
rect 1452 4604 1458 4616
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1452 4576 1593 4604
rect 1452 4564 1458 4576
rect 1581 4573 1593 4576
rect 1627 4573 1639 4607
rect 3970 4604 3976 4616
rect 3931 4576 3976 4604
rect 1581 4567 1639 4573
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4617 4607 4675 4613
rect 4617 4573 4629 4607
rect 4663 4573 4675 4607
rect 5902 4604 5908 4616
rect 5863 4576 5908 4604
rect 4617 4567 4675 4573
rect 4632 4536 4660 4567
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 8202 4564 8208 4616
rect 8260 4604 8266 4616
rect 9401 4607 9459 4613
rect 9401 4604 9413 4607
rect 8260 4576 9413 4604
rect 8260 4564 8266 4576
rect 9401 4573 9413 4576
rect 9447 4573 9459 4607
rect 9858 4604 9864 4616
rect 9819 4576 9864 4604
rect 9401 4567 9459 4573
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 15194 4604 15200 4616
rect 15155 4576 15200 4604
rect 15194 4564 15200 4576
rect 15252 4564 15258 4616
rect 22373 4607 22431 4613
rect 22373 4573 22385 4607
rect 22419 4604 22431 4607
rect 24394 4604 24400 4616
rect 22419 4576 24400 4604
rect 22419 4573 22431 4576
rect 22373 4567 22431 4573
rect 24394 4564 24400 4576
rect 24452 4564 24458 4616
rect 34885 4607 34943 4613
rect 34885 4573 34897 4607
rect 34931 4604 34943 4607
rect 35345 4607 35403 4613
rect 35345 4604 35357 4607
rect 34931 4576 35357 4604
rect 34931 4573 34943 4576
rect 34885 4567 34943 4573
rect 35345 4573 35357 4576
rect 35391 4573 35403 4607
rect 35345 4567 35403 4573
rect 37366 4564 37372 4616
rect 37424 4604 37430 4616
rect 37645 4607 37703 4613
rect 37645 4604 37657 4607
rect 37424 4576 37657 4604
rect 37424 4564 37430 4576
rect 37645 4573 37657 4576
rect 37691 4573 37703 4607
rect 37645 4567 37703 4573
rect 5810 4536 5816 4548
rect 4632 4508 5816 4536
rect 5810 4496 5816 4508
rect 5868 4496 5874 4548
rect 6549 4539 6607 4545
rect 6549 4505 6561 4539
rect 6595 4536 6607 4539
rect 7282 4536 7288 4548
rect 6595 4508 7288 4536
rect 6595 4505 6607 4508
rect 6549 4499 6607 4505
rect 7282 4496 7288 4508
rect 7340 4496 7346 4548
rect 15378 4536 15384 4548
rect 15339 4508 15384 4536
rect 15378 4496 15384 4508
rect 15436 4496 15442 4548
rect 9306 4468 9312 4480
rect 9267 4440 9312 4468
rect 9306 4428 9312 4440
rect 9364 4428 9370 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 3970 4224 3976 4276
rect 4028 4264 4034 4276
rect 4028 4236 13124 4264
rect 4028 4224 4034 4236
rect 9490 4196 9496 4208
rect 7392 4168 9496 4196
rect 7392 4140 7420 4168
rect 9490 4156 9496 4168
rect 9548 4156 9554 4208
rect 13096 4196 13124 4236
rect 15378 4224 15384 4276
rect 15436 4264 15442 4276
rect 15565 4267 15623 4273
rect 15565 4264 15577 4267
rect 15436 4236 15577 4264
rect 15436 4224 15442 4236
rect 15565 4233 15577 4236
rect 15611 4233 15623 4267
rect 15565 4227 15623 4233
rect 15746 4196 15752 4208
rect 11624 4168 11836 4196
rect 13096 4168 15752 4196
rect 4706 4128 4712 4140
rect 4667 4100 4712 4128
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 6549 4131 6607 4137
rect 6549 4097 6561 4131
rect 6595 4128 6607 4131
rect 7098 4128 7104 4140
rect 6595 4100 7104 4128
rect 6595 4097 6607 4100
rect 6549 4091 6607 4097
rect 7098 4088 7104 4100
rect 7156 4088 7162 4140
rect 7282 4128 7288 4140
rect 7243 4100 7288 4128
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 7432 4100 7477 4128
rect 7432 4088 7438 4100
rect 1946 4060 1952 4072
rect 1907 4032 1952 4060
rect 1946 4020 1952 4032
rect 2004 4020 2010 4072
rect 2133 4063 2191 4069
rect 2133 4029 2145 4063
rect 2179 4060 2191 4063
rect 2498 4060 2504 4072
rect 2179 4032 2504 4060
rect 2179 4029 2191 4032
rect 2133 4023 2191 4029
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 2593 4063 2651 4069
rect 2593 4029 2605 4063
rect 2639 4029 2651 4063
rect 2593 4023 2651 4029
rect 8021 4063 8079 4069
rect 8021 4029 8033 4063
rect 8067 4060 8079 4063
rect 8481 4063 8539 4069
rect 8481 4060 8493 4063
rect 8067 4032 8493 4060
rect 8067 4029 8079 4032
rect 8021 4023 8079 4029
rect 8481 4029 8493 4032
rect 8527 4029 8539 4063
rect 8662 4060 8668 4072
rect 8623 4032 8668 4060
rect 8481 4023 8539 4029
rect 658 3952 664 4004
rect 716 3992 722 4004
rect 2608 3992 2636 4023
rect 8662 4020 8668 4032
rect 8720 4020 8726 4072
rect 9309 4063 9367 4069
rect 9309 4060 9321 4063
rect 9232 4032 9321 4060
rect 716 3964 2636 3992
rect 716 3952 722 3964
rect 4798 3924 4804 3936
rect 4759 3896 4804 3924
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 5350 3924 5356 3936
rect 5311 3896 5356 3924
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 6546 3924 6552 3936
rect 6503 3896 6552 3924
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 6638 3884 6644 3936
rect 6696 3924 6702 3936
rect 9232 3924 9260 4032
rect 9309 4029 9321 4032
rect 9355 4029 9367 4063
rect 9309 4023 9367 4029
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 11624 4060 11652 4168
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4097 11759 4131
rect 11701 4091 11759 4097
rect 9456 4032 11652 4060
rect 9456 4020 9462 4032
rect 9490 3952 9496 4004
rect 9548 3992 9554 4004
rect 11716 3992 11744 4091
rect 11808 4060 11836 4168
rect 15746 4156 15752 4168
rect 15804 4196 15810 4208
rect 23658 4196 23664 4208
rect 15804 4168 23664 4196
rect 15804 4156 15810 4168
rect 23658 4156 23664 4168
rect 23716 4156 23722 4208
rect 34808 4168 36216 4196
rect 15654 4128 15660 4140
rect 15615 4100 15660 4128
rect 15654 4088 15660 4100
rect 15712 4088 15718 4140
rect 20346 4128 20352 4140
rect 20307 4100 20352 4128
rect 20346 4088 20352 4100
rect 20404 4088 20410 4140
rect 22186 4128 22192 4140
rect 21652 4100 22192 4128
rect 21652 4060 21680 4100
rect 22186 4088 22192 4100
rect 22244 4088 22250 4140
rect 32214 4128 32220 4140
rect 32175 4100 32220 4128
rect 32214 4088 32220 4100
rect 32272 4088 32278 4140
rect 34808 4128 34836 4168
rect 32508 4100 34836 4128
rect 36188 4128 36216 4168
rect 37274 4128 37280 4140
rect 36188 4100 37280 4128
rect 32508 4072 32536 4100
rect 37274 4088 37280 4100
rect 37332 4088 37338 4140
rect 37369 4131 37427 4137
rect 37369 4097 37381 4131
rect 37415 4097 37427 4131
rect 37369 4091 37427 4097
rect 11808 4032 21680 4060
rect 22554 4020 22560 4072
rect 22612 4060 22618 4072
rect 23385 4063 23443 4069
rect 23385 4060 23397 4063
rect 22612 4032 23397 4060
rect 22612 4020 22618 4032
rect 23385 4029 23397 4032
rect 23431 4029 23443 4063
rect 23566 4060 23572 4072
rect 23527 4032 23572 4060
rect 23385 4023 23443 4029
rect 23566 4020 23572 4032
rect 23624 4020 23630 4072
rect 23842 4060 23848 4072
rect 23803 4032 23848 4060
rect 23842 4020 23848 4032
rect 23900 4020 23906 4072
rect 32490 4060 32496 4072
rect 32451 4032 32496 4060
rect 32490 4020 32496 4032
rect 32548 4020 32554 4072
rect 34146 4020 34152 4072
rect 34204 4060 34210 4072
rect 34793 4063 34851 4069
rect 34793 4060 34805 4063
rect 34204 4032 34805 4060
rect 34204 4020 34210 4032
rect 34793 4029 34805 4032
rect 34839 4029 34851 4063
rect 34974 4060 34980 4072
rect 34935 4032 34980 4060
rect 34793 4023 34851 4029
rect 34974 4020 34980 4032
rect 35032 4020 35038 4072
rect 35434 4060 35440 4072
rect 35395 4032 35440 4060
rect 35434 4020 35440 4032
rect 35492 4020 35498 4072
rect 9548 3964 11744 3992
rect 9548 3952 9554 3964
rect 13814 3952 13820 4004
rect 13872 3992 13878 4004
rect 14826 3992 14832 4004
rect 13872 3964 14832 3992
rect 13872 3952 13878 3964
rect 14826 3952 14832 3964
rect 14884 3992 14890 4004
rect 37384 3992 37412 4091
rect 14884 3964 37412 3992
rect 14884 3952 14890 3964
rect 6696 3896 9260 3924
rect 6696 3884 6702 3896
rect 10410 3884 10416 3936
rect 10468 3924 10474 3936
rect 10781 3927 10839 3933
rect 10781 3924 10793 3927
rect 10468 3896 10793 3924
rect 10468 3884 10474 3896
rect 10781 3893 10793 3896
rect 10827 3893 10839 3927
rect 10781 3887 10839 3893
rect 11793 3927 11851 3933
rect 11793 3893 11805 3927
rect 11839 3924 11851 3927
rect 11882 3924 11888 3936
rect 11839 3896 11888 3924
rect 11839 3893 11851 3896
rect 11793 3887 11851 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 18138 3924 18144 3936
rect 18099 3896 18144 3924
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 20162 3884 20168 3936
rect 20220 3924 20226 3936
rect 20257 3927 20315 3933
rect 20257 3924 20269 3927
rect 20220 3896 20269 3924
rect 20220 3884 20226 3896
rect 20257 3893 20269 3896
rect 20303 3893 20315 3927
rect 20257 3887 20315 3893
rect 22281 3927 22339 3933
rect 22281 3893 22293 3927
rect 22327 3924 22339 3927
rect 24578 3924 24584 3936
rect 22327 3896 24584 3924
rect 22327 3893 22339 3896
rect 22281 3887 22339 3893
rect 24578 3884 24584 3896
rect 24636 3884 24642 3936
rect 37274 3884 37280 3936
rect 37332 3924 37338 3936
rect 37461 3927 37519 3933
rect 37461 3924 37473 3927
rect 37332 3896 37473 3924
rect 37332 3884 37338 3896
rect 37461 3893 37473 3896
rect 37507 3893 37519 3927
rect 37461 3887 37519 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 2498 3720 2504 3732
rect 2459 3692 2504 3720
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 3068 3692 5488 3720
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3516 2007 3519
rect 2130 3516 2136 3528
rect 1995 3488 2136 3516
rect 1995 3485 2007 3488
rect 1949 3479 2007 3485
rect 2130 3476 2136 3488
rect 2188 3476 2194 3528
rect 3068 3525 3096 3692
rect 5350 3652 5356 3664
rect 4632 3624 5356 3652
rect 4632 3593 4660 3624
rect 5350 3612 5356 3624
rect 5408 3612 5414 3664
rect 5460 3652 5488 3692
rect 8662 3680 8668 3732
rect 8720 3720 8726 3732
rect 9217 3723 9275 3729
rect 9217 3720 9229 3723
rect 8720 3692 9229 3720
rect 8720 3680 8726 3692
rect 9217 3689 9229 3692
rect 9263 3689 9275 3723
rect 32490 3720 32496 3732
rect 9217 3683 9275 3689
rect 12406 3692 32496 3720
rect 12406 3652 12434 3692
rect 32490 3680 32496 3692
rect 32548 3680 32554 3732
rect 34146 3720 34152 3732
rect 34107 3692 34152 3720
rect 34146 3680 34152 3692
rect 34204 3680 34210 3732
rect 34790 3680 34796 3732
rect 34848 3720 34854 3732
rect 35069 3723 35127 3729
rect 35069 3720 35081 3723
rect 34848 3692 35081 3720
rect 34848 3680 34854 3692
rect 35069 3689 35081 3692
rect 35115 3689 35127 3723
rect 35069 3683 35127 3689
rect 5460 3624 12434 3652
rect 15105 3655 15163 3661
rect 15105 3621 15117 3655
rect 15151 3652 15163 3655
rect 15194 3652 15200 3664
rect 15151 3624 15200 3652
rect 15151 3621 15163 3624
rect 15105 3615 15163 3621
rect 15194 3612 15200 3624
rect 15252 3612 15258 3664
rect 22554 3652 22560 3664
rect 16546 3624 18736 3652
rect 22515 3624 22560 3652
rect 4617 3587 4675 3593
rect 4617 3553 4629 3587
rect 4663 3553 4675 3587
rect 4798 3584 4804 3596
rect 4759 3556 4804 3584
rect 4617 3547 4675 3553
rect 4798 3544 4804 3556
rect 4856 3544 4862 3596
rect 5166 3584 5172 3596
rect 5127 3556 5172 3584
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 10226 3584 10232 3596
rect 8312 3556 10232 3584
rect 2593 3519 2651 3525
rect 2593 3485 2605 3519
rect 2639 3516 2651 3519
rect 3053 3519 3111 3525
rect 3053 3516 3065 3519
rect 2639 3488 3065 3516
rect 2639 3485 2651 3488
rect 2593 3479 2651 3485
rect 3053 3485 3065 3488
rect 3099 3485 3111 3519
rect 3053 3479 3111 3485
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 2958 3408 2964 3460
rect 3016 3448 3022 3460
rect 3804 3448 3832 3479
rect 7006 3476 7012 3528
rect 7064 3516 7070 3528
rect 8312 3525 8340 3556
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 10410 3584 10416 3596
rect 10371 3556 10416 3584
rect 10410 3544 10416 3556
rect 10468 3544 10474 3596
rect 10962 3584 10968 3596
rect 10923 3556 10968 3584
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 16546 3584 16574 3624
rect 16758 3584 16764 3596
rect 12406 3556 16574 3584
rect 16719 3556 16764 3584
rect 7101 3519 7159 3525
rect 7101 3516 7113 3519
rect 7064 3488 7113 3516
rect 7064 3476 7070 3488
rect 7101 3485 7113 3488
rect 7147 3485 7159 3519
rect 7101 3479 7159 3485
rect 8297 3519 8355 3525
rect 8297 3485 8309 3519
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9766 3516 9772 3528
rect 9355 3488 9772 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 3016 3420 3832 3448
rect 7116 3448 7144 3479
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 9861 3451 9919 3457
rect 7116 3420 9812 3448
rect 3016 3408 3022 3420
rect 1578 3340 1584 3392
rect 1636 3380 1642 3392
rect 1857 3383 1915 3389
rect 1857 3380 1869 3383
rect 1636 3352 1869 3380
rect 1636 3340 1642 3352
rect 1857 3349 1869 3352
rect 1903 3349 1915 3383
rect 3142 3380 3148 3392
rect 3103 3352 3148 3380
rect 1857 3343 1915 3349
rect 3142 3340 3148 3352
rect 3200 3340 3206 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 7009 3383 7067 3389
rect 7009 3380 7021 3383
rect 6880 3352 7021 3380
rect 6880 3340 6886 3352
rect 7009 3349 7021 3352
rect 7055 3349 7067 3383
rect 7009 3343 7067 3349
rect 8205 3383 8263 3389
rect 8205 3349 8217 3383
rect 8251 3380 8263 3383
rect 9122 3380 9128 3392
rect 8251 3352 9128 3380
rect 8251 3349 8263 3352
rect 8205 3343 8263 3349
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 9784 3380 9812 3420
rect 9861 3417 9873 3451
rect 9907 3448 9919 3451
rect 10597 3451 10655 3457
rect 10597 3448 10609 3451
rect 9907 3420 10609 3448
rect 9907 3417 9919 3420
rect 9861 3411 9919 3417
rect 10597 3417 10609 3420
rect 10643 3417 10655 3451
rect 12406 3448 12434 3556
rect 16758 3544 16764 3556
rect 16816 3544 16822 3596
rect 12713 3519 12771 3525
rect 12713 3485 12725 3519
rect 12759 3485 12771 3519
rect 15562 3516 15568 3528
rect 15523 3488 15568 3516
rect 12713 3479 12771 3485
rect 10597 3411 10655 3417
rect 11624 3420 12434 3448
rect 11624 3380 11652 3420
rect 9784 3352 11652 3380
rect 11698 3340 11704 3392
rect 11756 3380 11762 3392
rect 12728 3380 12756 3479
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 16206 3516 16212 3528
rect 16167 3488 16212 3516
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 18708 3525 18736 3624
rect 22554 3612 22560 3624
rect 22612 3612 22618 3664
rect 23109 3655 23167 3661
rect 23109 3621 23121 3655
rect 23155 3652 23167 3655
rect 23566 3652 23572 3664
rect 23155 3624 23572 3652
rect 23155 3621 23167 3624
rect 23109 3615 23167 3621
rect 23566 3612 23572 3624
rect 23624 3612 23630 3664
rect 23676 3624 24900 3652
rect 20162 3584 20168 3596
rect 20123 3556 20168 3584
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 20622 3584 20628 3596
rect 20583 3556 20628 3584
rect 20622 3544 20628 3556
rect 20680 3544 20686 3596
rect 23676 3584 23704 3624
rect 24394 3584 24400 3596
rect 22572 3556 23704 3584
rect 24355 3556 24400 3584
rect 22572 3528 22600 3556
rect 24394 3544 24400 3556
rect 24452 3544 24458 3596
rect 24578 3584 24584 3596
rect 24539 3556 24584 3584
rect 24578 3544 24584 3556
rect 24636 3544 24642 3596
rect 24872 3593 24900 3624
rect 24857 3587 24915 3593
rect 24857 3553 24869 3587
rect 24903 3553 24915 3587
rect 32214 3584 32220 3596
rect 24857 3547 24915 3553
rect 25792 3556 32220 3584
rect 18693 3519 18751 3525
rect 18693 3485 18705 3519
rect 18739 3516 18751 3519
rect 18782 3516 18788 3528
rect 18739 3488 18788 3516
rect 18739 3485 18751 3488
rect 18693 3479 18751 3485
rect 18782 3476 18788 3488
rect 18840 3476 18846 3528
rect 19521 3519 19579 3525
rect 19521 3485 19533 3519
rect 19567 3516 19579 3519
rect 19981 3519 20039 3525
rect 19981 3516 19993 3519
rect 19567 3488 19993 3516
rect 19567 3485 19579 3488
rect 19521 3479 19579 3485
rect 19981 3485 19993 3488
rect 20027 3485 20039 3519
rect 19981 3479 20039 3485
rect 22554 3476 22560 3528
rect 22612 3476 22618 3528
rect 23014 3516 23020 3528
rect 22975 3488 23020 3516
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 23658 3516 23664 3528
rect 23619 3488 23664 3516
rect 23658 3476 23664 3488
rect 23716 3516 23722 3528
rect 24118 3516 24124 3528
rect 23716 3488 24124 3516
rect 23716 3476 23722 3488
rect 24118 3476 24124 3488
rect 24176 3476 24182 3528
rect 15657 3451 15715 3457
rect 15657 3417 15669 3451
rect 15703 3448 15715 3451
rect 16393 3451 16451 3457
rect 16393 3448 16405 3451
rect 15703 3420 16405 3448
rect 15703 3417 15715 3420
rect 15657 3411 15715 3417
rect 16393 3417 16405 3420
rect 16439 3417 16451 3451
rect 23032 3448 23060 3476
rect 25792 3448 25820 3556
rect 32214 3544 32220 3556
rect 32272 3544 32278 3596
rect 37458 3584 37464 3596
rect 35176 3556 37464 3584
rect 28169 3519 28227 3525
rect 28169 3516 28181 3519
rect 23032 3420 25820 3448
rect 26206 3488 28181 3516
rect 16393 3411 16451 3417
rect 11756 3352 12756 3380
rect 11756 3340 11762 3352
rect 18322 3340 18328 3392
rect 18380 3380 18386 3392
rect 18601 3383 18659 3389
rect 18601 3380 18613 3383
rect 18380 3352 18613 3380
rect 18380 3340 18386 3352
rect 18601 3349 18613 3352
rect 18647 3349 18659 3383
rect 18601 3343 18659 3349
rect 23753 3383 23811 3389
rect 23753 3349 23765 3383
rect 23799 3380 23811 3383
rect 24026 3380 24032 3392
rect 23799 3352 24032 3380
rect 23799 3349 23811 3352
rect 23753 3343 23811 3349
rect 24026 3340 24032 3352
rect 24084 3340 24090 3392
rect 24118 3340 24124 3392
rect 24176 3380 24182 3392
rect 26206 3380 26234 3488
rect 28169 3485 28181 3488
rect 28215 3485 28227 3519
rect 28169 3479 28227 3485
rect 28629 3519 28687 3525
rect 28629 3485 28641 3519
rect 28675 3485 28687 3519
rect 28629 3479 28687 3485
rect 27798 3408 27804 3460
rect 27856 3448 27862 3460
rect 28644 3448 28672 3479
rect 32582 3476 32588 3528
rect 32640 3516 32646 3528
rect 32677 3519 32735 3525
rect 32677 3516 32689 3519
rect 32640 3488 32689 3516
rect 32640 3476 32646 3488
rect 32677 3485 32689 3488
rect 32723 3485 32735 3519
rect 32677 3479 32735 3485
rect 33226 3476 33232 3528
rect 33284 3516 33290 3528
rect 35176 3525 35204 3556
rect 37458 3544 37464 3556
rect 37516 3544 37522 3596
rect 33321 3519 33379 3525
rect 33321 3516 33333 3519
rect 33284 3488 33333 3516
rect 33284 3476 33290 3488
rect 33321 3485 33333 3488
rect 33367 3485 33379 3519
rect 33321 3479 33379 3485
rect 35161 3519 35219 3525
rect 35161 3485 35173 3519
rect 35207 3485 35219 3519
rect 35618 3516 35624 3528
rect 35579 3488 35624 3516
rect 35161 3479 35219 3485
rect 35618 3476 35624 3488
rect 35676 3476 35682 3528
rect 38102 3476 38108 3528
rect 38160 3516 38166 3528
rect 38160 3488 38205 3516
rect 38160 3476 38166 3488
rect 27856 3420 28672 3448
rect 27856 3408 27862 3420
rect 35802 3408 35808 3460
rect 35860 3448 35866 3460
rect 36265 3451 36323 3457
rect 36265 3448 36277 3451
rect 35860 3420 36277 3448
rect 35860 3408 35866 3420
rect 36265 3417 36277 3420
rect 36311 3417 36323 3451
rect 36265 3411 36323 3417
rect 37458 3408 37464 3460
rect 37516 3448 37522 3460
rect 37921 3451 37979 3457
rect 37921 3448 37933 3451
rect 37516 3420 37933 3448
rect 37516 3408 37522 3420
rect 37921 3417 37933 3420
rect 37967 3417 37979 3451
rect 37921 3411 37979 3417
rect 24176 3352 26234 3380
rect 24176 3340 24182 3352
rect 27982 3340 27988 3392
rect 28040 3380 28046 3392
rect 28077 3383 28135 3389
rect 28077 3380 28089 3383
rect 28040 3352 28089 3380
rect 28040 3340 28046 3352
rect 28077 3349 28089 3352
rect 28123 3349 28135 3383
rect 28077 3343 28135 3349
rect 32769 3383 32827 3389
rect 32769 3349 32781 3383
rect 32815 3380 32827 3383
rect 33410 3380 33416 3392
rect 32815 3352 33416 3380
rect 32815 3349 32827 3352
rect 32769 3343 32827 3349
rect 33410 3340 33416 3352
rect 33468 3340 33474 3392
rect 35710 3380 35716 3392
rect 35671 3352 35716 3380
rect 35710 3340 35716 3352
rect 35768 3340 35774 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 5460 3148 6960 3176
rect 3142 3108 3148 3120
rect 3103 3080 3148 3108
rect 3142 3068 3148 3080
rect 3200 3068 3206 3120
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 2958 3040 2964 3052
rect 2919 3012 2964 3040
rect 2958 3000 2964 3012
rect 3016 3000 3022 3052
rect 5460 3049 5488 3148
rect 6822 3108 6828 3120
rect 6783 3080 6828 3108
rect 6822 3068 6828 3080
rect 6880 3068 6886 3120
rect 6932 3108 6960 3148
rect 7098 3136 7104 3188
rect 7156 3176 7162 3188
rect 13814 3176 13820 3188
rect 7156 3148 13820 3176
rect 7156 3136 7162 3148
rect 13814 3136 13820 3148
rect 13872 3136 13878 3188
rect 15654 3136 15660 3188
rect 15712 3176 15718 3188
rect 15712 3148 33548 3176
rect 15712 3136 15718 3148
rect 8294 3108 8300 3120
rect 6932 3080 8300 3108
rect 8294 3068 8300 3080
rect 8352 3068 8358 3120
rect 9122 3108 9128 3120
rect 9083 3080 9128 3108
rect 9122 3068 9128 3080
rect 9180 3068 9186 3120
rect 11882 3108 11888 3120
rect 11843 3080 11888 3108
rect 11882 3068 11888 3080
rect 11940 3068 11946 3120
rect 18322 3108 18328 3120
rect 18283 3080 18328 3108
rect 18322 3068 18328 3080
rect 18380 3068 18386 3120
rect 24026 3108 24032 3120
rect 23987 3080 24032 3108
rect 24026 3068 24032 3080
rect 24084 3068 24090 3120
rect 27982 3108 27988 3120
rect 27943 3080 27988 3108
rect 27982 3068 27988 3080
rect 28040 3068 28046 3120
rect 33410 3108 33416 3120
rect 33371 3080 33416 3108
rect 33410 3068 33416 3080
rect 33468 3068 33474 3120
rect 33520 3108 33548 3148
rect 35342 3136 35348 3188
rect 35400 3176 35406 3188
rect 36630 3176 36636 3188
rect 35400 3148 36636 3176
rect 35400 3136 35406 3148
rect 36630 3136 36636 3148
rect 36688 3136 36694 3188
rect 37458 3176 37464 3188
rect 37419 3148 37464 3176
rect 37458 3136 37464 3148
rect 37516 3136 37522 3188
rect 37550 3108 37556 3120
rect 33520 3080 37556 3108
rect 37550 3068 37556 3080
rect 37608 3068 37614 3120
rect 5445 3043 5503 3049
rect 5445 3009 5457 3043
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5902 3000 5908 3052
rect 5960 3040 5966 3052
rect 6641 3043 6699 3049
rect 6641 3040 6653 3043
rect 5960 3012 6653 3040
rect 5960 3000 5966 3012
rect 6641 3009 6653 3012
rect 6687 3009 6699 3043
rect 8938 3040 8944 3052
rect 8899 3012 8944 3040
rect 6641 3003 6699 3009
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 11698 3040 11704 3052
rect 11659 3012 11704 3040
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 16206 3000 16212 3052
rect 16264 3040 16270 3052
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16264 3012 16681 3040
rect 16264 3000 16270 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 18138 3040 18144 3052
rect 18099 3012 18144 3040
rect 16669 3003 16727 3009
rect 18138 3000 18144 3012
rect 18196 3000 18202 3052
rect 27798 3040 27804 3052
rect 27759 3012 27804 3040
rect 27798 3000 27804 3012
rect 27856 3000 27862 3052
rect 33226 3040 33232 3052
rect 33187 3012 33232 3040
rect 33226 3000 33232 3012
rect 33284 3000 33290 3052
rect 37369 3043 37427 3049
rect 37369 3009 37381 3043
rect 37415 3040 37427 3043
rect 37642 3040 37648 3052
rect 37415 3012 37648 3040
rect 37415 3009 37427 3012
rect 37369 3003 37427 3009
rect 37642 3000 37648 3012
rect 37700 3000 37706 3052
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 3421 2975 3479 2981
rect 3421 2972 3433 2975
rect 3292 2944 3433 2972
rect 3292 2932 3298 2944
rect 3421 2941 3433 2944
rect 3467 2941 3479 2975
rect 7098 2972 7104 2984
rect 7059 2944 7104 2972
rect 3421 2935 3479 2941
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 9401 2975 9459 2981
rect 9401 2941 9413 2975
rect 9447 2941 9459 2975
rect 12250 2972 12256 2984
rect 12211 2944 12256 2972
rect 9401 2935 9459 2941
rect 6454 2864 6460 2916
rect 6512 2904 6518 2916
rect 9416 2904 9444 2935
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 18690 2972 18696 2984
rect 18651 2944 18696 2972
rect 18690 2932 18696 2944
rect 18748 2932 18754 2984
rect 23385 2975 23443 2981
rect 23385 2941 23397 2975
rect 23431 2972 23443 2975
rect 23845 2975 23903 2981
rect 23845 2972 23857 2975
rect 23431 2944 23857 2972
rect 23431 2941 23443 2944
rect 23385 2935 23443 2941
rect 23845 2941 23857 2944
rect 23891 2941 23903 2975
rect 24486 2972 24492 2984
rect 24447 2944 24492 2972
rect 23845 2935 23903 2941
rect 24486 2932 24492 2944
rect 24544 2932 24550 2984
rect 28350 2972 28356 2984
rect 24596 2944 26234 2972
rect 28311 2944 28356 2972
rect 6512 2876 9444 2904
rect 6512 2864 6518 2876
rect 18782 2864 18788 2916
rect 18840 2904 18846 2916
rect 24596 2904 24624 2944
rect 18840 2876 24624 2904
rect 26206 2904 26234 2944
rect 28350 2932 28356 2944
rect 28408 2932 28414 2984
rect 35069 2975 35127 2981
rect 35069 2941 35081 2975
rect 35115 2972 35127 2975
rect 35526 2972 35532 2984
rect 35115 2944 35532 2972
rect 35115 2941 35127 2944
rect 35069 2935 35127 2941
rect 35526 2932 35532 2944
rect 35584 2932 35590 2984
rect 32582 2904 32588 2916
rect 26206 2876 32588 2904
rect 18840 2864 18846 2876
rect 32582 2864 32588 2876
rect 32640 2864 32646 2916
rect 5353 2839 5411 2845
rect 5353 2805 5365 2839
rect 5399 2836 5411 2839
rect 5626 2836 5632 2848
rect 5399 2808 5632 2836
rect 5399 2805 5411 2808
rect 5353 2799 5411 2805
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 22186 2796 22192 2848
rect 22244 2836 22250 2848
rect 32674 2836 32680 2848
rect 22244 2808 32680 2836
rect 22244 2796 22250 2808
rect 32674 2796 32680 2808
rect 32732 2796 32738 2848
rect 33686 2796 33692 2848
rect 33744 2836 33750 2848
rect 35342 2836 35348 2848
rect 33744 2808 35348 2836
rect 33744 2796 33750 2808
rect 35342 2796 35348 2808
rect 35400 2796 35406 2848
rect 35986 2836 35992 2848
rect 35947 2808 35992 2836
rect 35986 2796 35992 2808
rect 36044 2796 36050 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 21726 2592 21732 2644
rect 21784 2632 21790 2644
rect 22005 2635 22063 2641
rect 22005 2632 22017 2635
rect 21784 2604 22017 2632
rect 21784 2592 21790 2604
rect 22005 2601 22017 2604
rect 22051 2601 22063 2635
rect 22005 2595 22063 2601
rect 37829 2635 37887 2641
rect 37829 2601 37841 2635
rect 37875 2632 37887 2635
rect 38102 2632 38108 2644
rect 37875 2604 38108 2632
rect 37875 2601 37887 2604
rect 37829 2595 37887 2601
rect 38102 2592 38108 2604
rect 38160 2592 38166 2644
rect 4522 2524 4528 2576
rect 4580 2564 4586 2576
rect 9858 2564 9864 2576
rect 4580 2536 6868 2564
rect 4580 2524 4586 2536
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 1578 2496 1584 2508
rect 1539 2468 1584 2496
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 2774 2496 2780 2508
rect 2735 2468 2780 2496
rect 2774 2456 2780 2468
rect 2832 2456 2838 2508
rect 5626 2496 5632 2508
rect 5587 2468 5632 2496
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 5810 2496 5816 2508
rect 5771 2468 5816 2496
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 6178 2456 6184 2508
rect 6236 2496 6242 2508
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 6236 2468 6377 2496
rect 6236 2456 6242 2468
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6546 2496 6552 2508
rect 6507 2468 6552 2496
rect 6365 2459 6423 2465
rect 6546 2456 6552 2468
rect 6604 2456 6610 2508
rect 6840 2505 6868 2536
rect 9048 2536 9864 2564
rect 9048 2505 9076 2536
rect 9858 2524 9864 2536
rect 9916 2524 9922 2576
rect 37366 2564 37372 2576
rect 34164 2536 37372 2564
rect 6825 2499 6883 2505
rect 6825 2465 6837 2499
rect 6871 2465 6883 2499
rect 6825 2459 6883 2465
rect 9033 2499 9091 2505
rect 9033 2465 9045 2499
rect 9079 2465 9091 2499
rect 9033 2459 9091 2465
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 9306 2496 9312 2508
rect 9263 2468 9312 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 9674 2496 9680 2508
rect 9635 2468 9680 2496
rect 9674 2456 9680 2468
rect 9732 2456 9738 2508
rect 33686 2496 33692 2508
rect 33647 2468 33692 2496
rect 33686 2456 33692 2468
rect 33744 2456 33750 2508
rect 34164 2505 34192 2536
rect 37366 2524 37372 2536
rect 37424 2524 37430 2576
rect 34149 2499 34207 2505
rect 34149 2465 34161 2499
rect 34195 2465 34207 2499
rect 34149 2459 34207 2465
rect 34885 2499 34943 2505
rect 34885 2465 34897 2499
rect 34931 2496 34943 2499
rect 35986 2496 35992 2508
rect 34931 2468 35992 2496
rect 34931 2465 34943 2468
rect 34885 2459 34943 2465
rect 35986 2456 35992 2468
rect 36044 2456 36050 2508
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 21324 2400 21833 2428
rect 21324 2388 21330 2400
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 3878 2320 3884 2372
rect 3936 2360 3942 2372
rect 3973 2363 4031 2369
rect 3973 2360 3985 2363
rect 3936 2332 3985 2360
rect 3936 2320 3942 2332
rect 3973 2329 3985 2332
rect 4019 2329 4031 2363
rect 3973 2323 4031 2329
rect 33965 2363 34023 2369
rect 33965 2329 33977 2363
rect 34011 2329 34023 2363
rect 33965 2323 34023 2329
rect 35069 2363 35127 2369
rect 35069 2329 35081 2363
rect 35115 2360 35127 2363
rect 35710 2360 35716 2372
rect 35115 2332 35716 2360
rect 35115 2329 35127 2332
rect 35069 2323 35127 2329
rect 33980 2292 34008 2323
rect 35710 2320 35716 2332
rect 35768 2320 35774 2372
rect 36722 2360 36728 2372
rect 36683 2332 36728 2360
rect 36722 2320 36728 2332
rect 36780 2320 36786 2372
rect 37274 2292 37280 2304
rect 33980 2264 37280 2292
rect 37274 2252 37280 2264
rect 37332 2252 37338 2304
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 35900 47404 35952 47456
rect 37188 47404 37240 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 3332 47132 3384 47184
rect 1400 47107 1452 47116
rect 1400 47073 1409 47107
rect 1409 47073 1443 47107
rect 1443 47073 1452 47107
rect 1400 47064 1452 47073
rect 2872 47064 2924 47116
rect 4896 47064 4948 47116
rect 5172 47107 5224 47116
rect 5172 47073 5181 47107
rect 5181 47073 5215 47107
rect 5215 47073 5224 47107
rect 5172 47064 5224 47073
rect 20812 47132 20864 47184
rect 7380 47064 7432 47116
rect 17408 47107 17460 47116
rect 17408 47073 17417 47107
rect 17417 47073 17451 47107
rect 17451 47073 17460 47107
rect 17408 47064 17460 47073
rect 29736 47064 29788 47116
rect 32312 47064 32364 47116
rect 36728 47064 36780 47116
rect 8944 47039 8996 47048
rect 8944 47005 8953 47039
rect 8953 47005 8987 47039
rect 8987 47005 8996 47039
rect 8944 46996 8996 47005
rect 9772 47039 9824 47048
rect 9772 47005 9781 47039
rect 9781 47005 9815 47039
rect 9815 47005 9824 47039
rect 9772 46996 9824 47005
rect 16856 47039 16908 47048
rect 16856 47005 16865 47039
rect 16865 47005 16899 47039
rect 16899 47005 16908 47039
rect 16856 46996 16908 47005
rect 20168 46996 20220 47048
rect 3056 46971 3108 46980
rect 3056 46937 3065 46971
rect 3065 46937 3099 46971
rect 3099 46937 3108 46971
rect 3056 46928 3108 46937
rect 4620 46928 4672 46980
rect 8208 46971 8260 46980
rect 8208 46937 8217 46971
rect 8217 46937 8251 46971
rect 8251 46937 8260 46971
rect 8208 46928 8260 46937
rect 17040 46971 17092 46980
rect 17040 46937 17049 46971
rect 17049 46937 17083 46971
rect 17083 46937 17092 46971
rect 17040 46928 17092 46937
rect 19984 46860 20036 46912
rect 22100 46996 22152 47048
rect 24400 47039 24452 47048
rect 24400 47005 24409 47039
rect 24409 47005 24443 47039
rect 24443 47005 24452 47039
rect 24400 46996 24452 47005
rect 27988 47039 28040 47048
rect 27988 47005 27997 47039
rect 27997 47005 28031 47039
rect 28031 47005 28040 47039
rect 27988 46996 28040 47005
rect 29552 47039 29604 47048
rect 29552 47005 29561 47039
rect 29561 47005 29595 47039
rect 29595 47005 29604 47039
rect 29552 46996 29604 47005
rect 32128 47039 32180 47048
rect 32128 47005 32137 47039
rect 32137 47005 32171 47039
rect 32171 47005 32180 47039
rect 32128 46996 32180 47005
rect 36452 47039 36504 47048
rect 36452 47005 36461 47039
rect 36461 47005 36495 47039
rect 36495 47005 36504 47039
rect 36452 46996 36504 47005
rect 37740 47039 37792 47048
rect 37740 47005 37749 47039
rect 37749 47005 37783 47039
rect 37783 47005 37792 47039
rect 37740 46996 37792 47005
rect 29276 46928 29328 46980
rect 32312 46971 32364 46980
rect 32312 46937 32321 46971
rect 32321 46937 32355 46971
rect 32355 46937 32364 46971
rect 32312 46928 32364 46937
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 8208 46656 8260 46708
rect 2596 46588 2648 46640
rect 8392 46588 8444 46640
rect 33232 46588 33284 46640
rect 35348 46588 35400 46640
rect 8116 46520 8168 46572
rect 9772 46563 9824 46572
rect 9772 46529 9781 46563
rect 9781 46529 9815 46563
rect 9815 46529 9824 46563
rect 9772 46520 9824 46529
rect 16856 46520 16908 46572
rect 20536 46563 20588 46572
rect 20536 46529 20545 46563
rect 20545 46529 20579 46563
rect 20579 46529 20588 46563
rect 20536 46520 20588 46529
rect 21180 46563 21232 46572
rect 21180 46529 21189 46563
rect 21189 46529 21223 46563
rect 21223 46529 21232 46563
rect 21180 46520 21232 46529
rect 22100 46563 22152 46572
rect 22100 46529 22109 46563
rect 22109 46529 22143 46563
rect 22143 46529 22152 46563
rect 22100 46520 22152 46529
rect 24400 46563 24452 46572
rect 24400 46529 24409 46563
rect 24409 46529 24443 46563
rect 24443 46529 24452 46563
rect 24400 46520 24452 46529
rect 27988 46563 28040 46572
rect 27988 46529 27997 46563
rect 27997 46529 28031 46563
rect 28031 46529 28040 46563
rect 27988 46520 28040 46529
rect 32128 46520 32180 46572
rect 36728 46563 36780 46572
rect 36728 46529 36737 46563
rect 36737 46529 36771 46563
rect 36771 46529 36780 46563
rect 36728 46520 36780 46529
rect 38016 46520 38068 46572
rect 2780 46452 2832 46504
rect 2964 46495 3016 46504
rect 2964 46461 2973 46495
rect 2973 46461 3007 46495
rect 3007 46461 3016 46495
rect 2964 46452 3016 46461
rect 5448 46452 5500 46504
rect 8208 46452 8260 46504
rect 18236 46495 18288 46504
rect 18236 46461 18245 46495
rect 18245 46461 18279 46495
rect 18279 46461 18288 46495
rect 18236 46452 18288 46461
rect 18696 46495 18748 46504
rect 18696 46461 18705 46495
rect 18705 46461 18739 46495
rect 18739 46461 18748 46495
rect 18696 46452 18748 46461
rect 22560 46452 22612 46504
rect 22652 46495 22704 46504
rect 22652 46461 22661 46495
rect 22661 46461 22695 46495
rect 22695 46461 22704 46495
rect 24584 46495 24636 46504
rect 22652 46452 22704 46461
rect 24584 46461 24593 46495
rect 24593 46461 24627 46495
rect 24627 46461 24636 46495
rect 24584 46452 24636 46461
rect 24492 46384 24544 46436
rect 28632 46452 28684 46504
rect 28356 46384 28408 46436
rect 33324 46452 33376 46504
rect 35808 46495 35860 46504
rect 35808 46461 35817 46495
rect 35817 46461 35851 46495
rect 35851 46461 35860 46495
rect 35808 46452 35860 46461
rect 33876 46384 33928 46436
rect 5816 46359 5868 46368
rect 5816 46325 5825 46359
rect 5825 46325 5859 46359
rect 5859 46325 5868 46359
rect 5816 46316 5868 46325
rect 6092 46316 6144 46368
rect 14924 46316 14976 46368
rect 19432 46316 19484 46368
rect 20352 46316 20404 46368
rect 21088 46316 21140 46368
rect 26240 46316 26292 46368
rect 30932 46359 30984 46368
rect 30932 46325 30941 46359
rect 30941 46325 30975 46359
rect 30975 46325 30984 46359
rect 30932 46316 30984 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 3056 46112 3108 46164
rect 4620 46155 4672 46164
rect 4620 46121 4629 46155
rect 4629 46121 4663 46155
rect 4663 46121 4672 46155
rect 4620 46112 4672 46121
rect 4896 46112 4948 46164
rect 8208 46155 8260 46164
rect 8208 46121 8217 46155
rect 8217 46121 8251 46155
rect 8251 46121 8260 46155
rect 8208 46112 8260 46121
rect 17040 46112 17092 46164
rect 18236 46155 18288 46164
rect 18236 46121 18245 46155
rect 18245 46121 18279 46155
rect 18279 46121 18288 46155
rect 18236 46112 18288 46121
rect 22560 46155 22612 46164
rect 22560 46121 22569 46155
rect 22569 46121 22603 46155
rect 22603 46121 22612 46155
rect 22560 46112 22612 46121
rect 24584 46112 24636 46164
rect 28632 46155 28684 46164
rect 28632 46121 28641 46155
rect 28641 46121 28675 46155
rect 28675 46121 28684 46155
rect 28632 46112 28684 46121
rect 29552 46155 29604 46164
rect 29552 46121 29561 46155
rect 29561 46121 29595 46155
rect 29595 46121 29604 46155
rect 29552 46112 29604 46121
rect 33324 46155 33376 46164
rect 33324 46121 33333 46155
rect 33333 46121 33367 46155
rect 33367 46121 33376 46155
rect 33324 46112 33376 46121
rect 33876 46155 33928 46164
rect 33876 46121 33885 46155
rect 33885 46121 33919 46155
rect 33919 46121 33928 46155
rect 33876 46112 33928 46121
rect 9036 46044 9088 46096
rect 20 45976 72 46028
rect 6092 45976 6144 46028
rect 6460 46019 6512 46028
rect 6460 45985 6469 46019
rect 6469 45985 6503 46019
rect 6503 45985 6512 46019
rect 6460 45976 6512 45985
rect 8944 46019 8996 46028
rect 8944 45985 8953 46019
rect 8953 45985 8987 46019
rect 8987 45985 8996 46019
rect 8944 45976 8996 45985
rect 14924 46019 14976 46028
rect 14924 45985 14933 46019
rect 14933 45985 14967 46019
rect 14967 45985 14976 46019
rect 14924 45976 14976 45985
rect 15476 46019 15528 46028
rect 15476 45985 15485 46019
rect 15485 45985 15519 46019
rect 15519 45985 15528 46019
rect 15476 45976 15528 45985
rect 20168 46019 20220 46028
rect 3240 45951 3292 45960
rect 3240 45917 3249 45951
rect 3249 45917 3283 45951
rect 3283 45917 3292 45951
rect 3240 45908 3292 45917
rect 4804 45908 4856 45960
rect 8116 45951 8168 45960
rect 8116 45917 8125 45951
rect 8125 45917 8159 45951
rect 8159 45917 8168 45951
rect 8116 45908 8168 45917
rect 17408 45951 17460 45960
rect 17408 45917 17417 45951
rect 17417 45917 17451 45951
rect 17451 45917 17460 45951
rect 17408 45908 17460 45917
rect 18052 45908 18104 45960
rect 20168 45985 20177 46019
rect 20177 45985 20211 46019
rect 20211 45985 20220 46019
rect 20168 45976 20220 45985
rect 20352 46019 20404 46028
rect 20352 45985 20361 46019
rect 20361 45985 20395 46019
rect 20395 45985 20404 46019
rect 20352 45976 20404 45985
rect 21272 46019 21324 46028
rect 21272 45985 21281 46019
rect 21281 45985 21315 46019
rect 21315 45985 21324 46019
rect 21272 45976 21324 45985
rect 26240 46019 26292 46028
rect 26240 45985 26249 46019
rect 26249 45985 26283 46019
rect 26283 45985 26292 46019
rect 27068 46019 27120 46028
rect 26240 45976 26292 45985
rect 27068 45985 27077 46019
rect 27077 45985 27111 46019
rect 27111 45985 27120 46019
rect 27068 45976 27120 45985
rect 30932 46019 30984 46028
rect 30932 45985 30941 46019
rect 30941 45985 30975 46019
rect 30975 45985 30984 46019
rect 30932 45976 30984 45985
rect 31576 45976 31628 46028
rect 36452 45976 36504 46028
rect 37372 46019 37424 46028
rect 37372 45985 37381 46019
rect 37381 45985 37415 46019
rect 37415 45985 37424 46019
rect 37372 45976 37424 45985
rect 22652 45951 22704 45960
rect 22652 45917 22661 45951
rect 22661 45917 22695 45951
rect 22695 45917 22704 45951
rect 22652 45908 22704 45917
rect 23848 45908 23900 45960
rect 28724 45951 28776 45960
rect 3056 45883 3108 45892
rect 3056 45849 3065 45883
rect 3065 45849 3099 45883
rect 3099 45849 3108 45883
rect 3056 45840 3108 45849
rect 5724 45840 5776 45892
rect 8944 45840 8996 45892
rect 15200 45840 15252 45892
rect 7472 45772 7524 45824
rect 8116 45772 8168 45824
rect 19340 45815 19392 45824
rect 19340 45781 19349 45815
rect 19349 45781 19383 45815
rect 19383 45781 19392 45815
rect 19340 45772 19392 45781
rect 28724 45917 28733 45951
rect 28733 45917 28767 45951
rect 28767 45917 28776 45951
rect 28724 45908 28776 45917
rect 33232 45951 33284 45960
rect 33232 45917 33241 45951
rect 33241 45917 33275 45951
rect 33275 45917 33284 45951
rect 33232 45908 33284 45917
rect 26424 45883 26476 45892
rect 26424 45849 26433 45883
rect 26433 45849 26467 45883
rect 26467 45849 26476 45883
rect 26424 45840 26476 45849
rect 31116 45883 31168 45892
rect 31116 45849 31125 45883
rect 31125 45849 31159 45883
rect 31159 45849 31168 45883
rect 31116 45840 31168 45849
rect 37372 45840 37424 45892
rect 38016 45772 38068 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 5724 45611 5776 45620
rect 5724 45577 5733 45611
rect 5733 45577 5767 45611
rect 5767 45577 5776 45611
rect 5724 45568 5776 45577
rect 8944 45611 8996 45620
rect 8944 45577 8953 45611
rect 8953 45577 8987 45611
rect 8987 45577 8996 45611
rect 8944 45568 8996 45577
rect 2780 45543 2832 45552
rect 2780 45509 2789 45543
rect 2789 45509 2823 45543
rect 2823 45509 2832 45543
rect 2780 45500 2832 45509
rect 2964 45432 3016 45484
rect 3240 45432 3292 45484
rect 6920 45500 6972 45552
rect 15200 45543 15252 45552
rect 15200 45509 15209 45543
rect 15209 45509 15243 45543
rect 15243 45509 15252 45543
rect 15200 45500 15252 45509
rect 19340 45500 19392 45552
rect 5816 45432 5868 45484
rect 8024 45432 8076 45484
rect 1400 45407 1452 45416
rect 1400 45373 1409 45407
rect 1409 45373 1443 45407
rect 1443 45373 1452 45407
rect 1400 45364 1452 45373
rect 1676 45407 1728 45416
rect 1676 45373 1685 45407
rect 1685 45373 1719 45407
rect 1719 45373 1728 45407
rect 1676 45364 1728 45373
rect 6736 45407 6788 45416
rect 6736 45373 6745 45407
rect 6745 45373 6779 45407
rect 6779 45373 6788 45407
rect 6736 45364 6788 45373
rect 8116 45407 8168 45416
rect 8116 45373 8125 45407
rect 8125 45373 8159 45407
rect 8159 45373 8168 45407
rect 8116 45364 8168 45373
rect 8852 45475 8904 45484
rect 8852 45441 8861 45475
rect 8861 45441 8895 45475
rect 8895 45441 8904 45475
rect 15292 45475 15344 45484
rect 8852 45432 8904 45441
rect 15292 45441 15301 45475
rect 15301 45441 15335 45475
rect 15335 45441 15344 45475
rect 15292 45432 15344 45441
rect 20076 45475 20128 45484
rect 20076 45441 20110 45475
rect 20110 45441 20128 45475
rect 20076 45432 20128 45441
rect 17960 45407 18012 45416
rect 2964 45296 3016 45348
rect 10048 45296 10100 45348
rect 17960 45373 17969 45407
rect 17969 45373 18003 45407
rect 18003 45373 18012 45407
rect 17960 45364 18012 45373
rect 19432 45364 19484 45416
rect 19800 45407 19852 45416
rect 19800 45373 19809 45407
rect 19809 45373 19843 45407
rect 19843 45373 19852 45407
rect 19800 45364 19852 45373
rect 22100 45432 22152 45484
rect 23020 45432 23072 45484
rect 20904 45228 20956 45280
rect 22192 45271 22244 45280
rect 22192 45237 22201 45271
rect 22201 45237 22235 45271
rect 22235 45237 22244 45271
rect 22192 45228 22244 45237
rect 22928 45296 22980 45348
rect 22836 45228 22888 45280
rect 26424 45568 26476 45620
rect 31116 45611 31168 45620
rect 31116 45577 31125 45611
rect 31125 45577 31159 45611
rect 31159 45577 31168 45611
rect 31116 45568 31168 45577
rect 29276 45543 29328 45552
rect 29276 45509 29285 45543
rect 29285 45509 29319 45543
rect 29319 45509 29328 45543
rect 29276 45500 29328 45509
rect 32312 45500 32364 45552
rect 37372 45543 37424 45552
rect 37372 45509 37381 45543
rect 37381 45509 37415 45543
rect 37415 45509 37424 45543
rect 37372 45500 37424 45509
rect 24768 45432 24820 45484
rect 24952 45432 25004 45484
rect 27160 45432 27212 45484
rect 31208 45432 31260 45484
rect 32404 45432 32456 45484
rect 37280 45475 37332 45484
rect 37280 45441 37289 45475
rect 37289 45441 37323 45475
rect 37323 45441 37332 45475
rect 37280 45432 37332 45441
rect 38384 45432 38436 45484
rect 28356 45407 28408 45416
rect 28356 45373 28365 45407
rect 28365 45373 28399 45407
rect 28399 45373 28408 45407
rect 28356 45364 28408 45373
rect 29276 45364 29328 45416
rect 35808 45407 35860 45416
rect 35808 45373 35817 45407
rect 35817 45373 35851 45407
rect 35851 45373 35860 45407
rect 35808 45364 35860 45373
rect 36544 45407 36596 45416
rect 36544 45373 36553 45407
rect 36553 45373 36587 45407
rect 36587 45373 36596 45407
rect 36544 45364 36596 45373
rect 36728 45407 36780 45416
rect 36728 45373 36737 45407
rect 36737 45373 36771 45407
rect 36771 45373 36780 45407
rect 36728 45364 36780 45373
rect 26884 45228 26936 45280
rect 37924 45228 37976 45280
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 2872 45024 2924 45076
rect 6736 45024 6788 45076
rect 7380 45067 7432 45076
rect 7380 45033 7389 45067
rect 7389 45033 7423 45067
rect 7423 45033 7432 45067
rect 7380 45024 7432 45033
rect 8852 45024 8904 45076
rect 37372 45024 37424 45076
rect 3056 44956 3108 45008
rect 23020 44956 23072 45008
rect 18144 44888 18196 44940
rect 19800 44888 19852 44940
rect 2504 44820 2556 44872
rect 6920 44820 6972 44872
rect 8208 44820 8260 44872
rect 19432 44820 19484 44872
rect 20720 44820 20772 44872
rect 2504 44684 2556 44736
rect 10508 44684 10560 44736
rect 19984 44684 20036 44736
rect 22376 44888 22428 44940
rect 27344 44956 27396 45008
rect 24768 44888 24820 44940
rect 37740 44956 37792 45008
rect 37096 44931 37148 44940
rect 37096 44897 37105 44931
rect 37105 44897 37139 44931
rect 37139 44897 37148 44931
rect 37096 44888 37148 44897
rect 37924 44931 37976 44940
rect 37924 44897 37933 44931
rect 37933 44897 37967 44931
rect 37967 44897 37976 44931
rect 37924 44888 37976 44897
rect 21088 44795 21140 44804
rect 21088 44761 21122 44795
rect 21122 44761 21140 44795
rect 21088 44752 21140 44761
rect 23572 44820 23624 44872
rect 22928 44795 22980 44804
rect 22100 44684 22152 44736
rect 22928 44761 22937 44795
rect 22937 44761 22971 44795
rect 22971 44761 22980 44795
rect 22928 44752 22980 44761
rect 23112 44752 23164 44804
rect 26056 44820 26108 44872
rect 24952 44752 25004 44804
rect 25780 44752 25832 44804
rect 22836 44727 22888 44736
rect 22836 44693 22845 44727
rect 22845 44693 22879 44727
rect 22879 44693 22888 44727
rect 22836 44684 22888 44693
rect 23020 44727 23072 44736
rect 23020 44693 23029 44727
rect 23029 44693 23063 44727
rect 23063 44693 23072 44727
rect 23020 44684 23072 44693
rect 23664 44727 23716 44736
rect 23664 44693 23673 44727
rect 23673 44693 23707 44727
rect 23707 44693 23716 44727
rect 23664 44684 23716 44693
rect 26976 44684 27028 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 20076 44480 20128 44532
rect 21180 44523 21232 44532
rect 21180 44489 21189 44523
rect 21189 44489 21223 44523
rect 21223 44489 21232 44523
rect 21180 44480 21232 44489
rect 23020 44480 23072 44532
rect 27160 44523 27212 44532
rect 27160 44489 27169 44523
rect 27169 44489 27203 44523
rect 27203 44489 27212 44523
rect 27160 44480 27212 44489
rect 36544 44480 36596 44532
rect 20720 44412 20772 44464
rect 18144 44387 18196 44396
rect 18144 44353 18153 44387
rect 18153 44353 18187 44387
rect 18187 44353 18196 44387
rect 18144 44344 18196 44353
rect 19248 44344 19300 44396
rect 19984 44387 20036 44396
rect 19984 44353 19993 44387
rect 19993 44353 20027 44387
rect 20027 44353 20036 44387
rect 19984 44344 20036 44353
rect 20904 44387 20956 44396
rect 20904 44353 20913 44387
rect 20913 44353 20947 44387
rect 20947 44353 20956 44387
rect 20904 44344 20956 44353
rect 23664 44412 23716 44464
rect 21456 44344 21508 44396
rect 23572 44387 23624 44396
rect 23572 44353 23581 44387
rect 23581 44353 23615 44387
rect 23615 44353 23624 44387
rect 23572 44344 23624 44353
rect 23940 44344 23992 44396
rect 24768 44344 24820 44396
rect 26056 44387 26108 44396
rect 26056 44353 26065 44387
rect 26065 44353 26099 44387
rect 26099 44353 26108 44387
rect 26056 44344 26108 44353
rect 26976 44387 27028 44396
rect 26976 44353 26985 44387
rect 26985 44353 27019 44387
rect 27019 44353 27028 44387
rect 26976 44344 27028 44353
rect 27804 44387 27856 44396
rect 27804 44353 27813 44387
rect 27813 44353 27847 44387
rect 27847 44353 27856 44387
rect 27804 44344 27856 44353
rect 29920 44387 29972 44396
rect 29920 44353 29929 44387
rect 29929 44353 29963 44387
rect 29963 44353 29972 44387
rect 29920 44344 29972 44353
rect 36728 44387 36780 44396
rect 36728 44353 36737 44387
rect 36737 44353 36771 44387
rect 36771 44353 36780 44387
rect 36728 44344 36780 44353
rect 37372 44387 37424 44396
rect 37372 44353 37381 44387
rect 37381 44353 37415 44387
rect 37415 44353 37424 44387
rect 37372 44344 37424 44353
rect 26240 44319 26292 44328
rect 26240 44285 26249 44319
rect 26249 44285 26283 44319
rect 26283 44285 26292 44319
rect 26240 44276 26292 44285
rect 29276 44208 29328 44260
rect 37372 44208 37424 44260
rect 19432 44140 19484 44192
rect 20260 44140 20312 44192
rect 25964 44140 26016 44192
rect 27988 44183 28040 44192
rect 27988 44149 27997 44183
rect 27997 44149 28031 44183
rect 28031 44149 28040 44183
rect 27988 44140 28040 44149
rect 29828 44140 29880 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 19248 43979 19300 43988
rect 19248 43945 19257 43979
rect 19257 43945 19291 43979
rect 19291 43945 19300 43979
rect 19248 43936 19300 43945
rect 23112 43936 23164 43988
rect 25780 43979 25832 43988
rect 25780 43945 25789 43979
rect 25789 43945 25823 43979
rect 25823 43945 25832 43979
rect 25780 43936 25832 43945
rect 27804 43936 27856 43988
rect 5448 43732 5500 43784
rect 22100 43800 22152 43852
rect 26056 43800 26108 43852
rect 38108 43843 38160 43852
rect 19432 43775 19484 43784
rect 19432 43741 19441 43775
rect 19441 43741 19475 43775
rect 19475 43741 19484 43775
rect 19432 43732 19484 43741
rect 21456 43732 21508 43784
rect 25780 43732 25832 43784
rect 25964 43775 26016 43784
rect 25964 43741 25973 43775
rect 25973 43741 26007 43775
rect 26007 43741 26016 43775
rect 25964 43732 26016 43741
rect 26884 43775 26936 43784
rect 26884 43741 26893 43775
rect 26893 43741 26927 43775
rect 26927 43741 26936 43775
rect 26884 43732 26936 43741
rect 38108 43809 38117 43843
rect 38117 43809 38151 43843
rect 38151 43809 38160 43843
rect 38108 43800 38160 43809
rect 27620 43775 27672 43784
rect 27620 43741 27629 43775
rect 27629 43741 27663 43775
rect 27663 43741 27672 43775
rect 27620 43732 27672 43741
rect 28356 43732 28408 43784
rect 29828 43775 29880 43784
rect 29828 43741 29862 43775
rect 29862 43741 29880 43775
rect 29828 43732 29880 43741
rect 36268 43775 36320 43784
rect 36268 43741 36277 43775
rect 36277 43741 36311 43775
rect 36311 43741 36320 43775
rect 36268 43732 36320 43741
rect 16672 43664 16724 43716
rect 27988 43664 28040 43716
rect 37464 43664 37516 43716
rect 17224 43639 17276 43648
rect 17224 43605 17233 43639
rect 17233 43605 17267 43639
rect 17267 43605 17276 43639
rect 17224 43596 17276 43605
rect 25136 43639 25188 43648
rect 25136 43605 25145 43639
rect 25145 43605 25179 43639
rect 25179 43605 25188 43639
rect 25136 43596 25188 43605
rect 29552 43596 29604 43648
rect 30932 43639 30984 43648
rect 30932 43605 30941 43639
rect 30941 43605 30975 43639
rect 30975 43605 30984 43639
rect 30932 43596 30984 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 19432 43435 19484 43444
rect 19432 43401 19441 43435
rect 19441 43401 19475 43435
rect 19475 43401 19484 43435
rect 19432 43392 19484 43401
rect 25780 43435 25832 43444
rect 25780 43401 25789 43435
rect 25789 43401 25823 43435
rect 25823 43401 25832 43435
rect 25780 43392 25832 43401
rect 26884 43392 26936 43444
rect 27344 43435 27396 43444
rect 27344 43401 27353 43435
rect 27353 43401 27387 43435
rect 27387 43401 27396 43435
rect 29920 43435 29972 43444
rect 27344 43392 27396 43401
rect 29920 43401 29929 43435
rect 29929 43401 29963 43435
rect 29963 43401 29972 43435
rect 29920 43392 29972 43401
rect 37464 43435 37516 43444
rect 37464 43401 37473 43435
rect 37473 43401 37507 43435
rect 37507 43401 37516 43435
rect 37464 43392 37516 43401
rect 17224 43324 17276 43376
rect 19984 43324 20036 43376
rect 20168 43299 20220 43308
rect 16580 43188 16632 43240
rect 20168 43265 20177 43299
rect 20177 43265 20211 43299
rect 20211 43265 20220 43299
rect 20168 43256 20220 43265
rect 23940 43299 23992 43308
rect 23940 43265 23949 43299
rect 23949 43265 23983 43299
rect 23983 43265 23992 43299
rect 23940 43256 23992 43265
rect 24032 43256 24084 43308
rect 26056 43324 26108 43376
rect 27068 43256 27120 43308
rect 29552 43299 29604 43308
rect 29552 43265 29561 43299
rect 29561 43265 29595 43299
rect 29595 43265 29604 43299
rect 29552 43256 29604 43265
rect 30288 43256 30340 43308
rect 31116 43299 31168 43308
rect 31116 43265 31125 43299
rect 31125 43265 31159 43299
rect 31159 43265 31168 43299
rect 31116 43256 31168 43265
rect 35808 43256 35860 43308
rect 36268 43256 36320 43308
rect 37832 43256 37884 43308
rect 20260 43188 20312 43240
rect 21180 43188 21232 43240
rect 21456 43120 21508 43172
rect 26240 43120 26292 43172
rect 26976 43163 27028 43172
rect 26976 43129 26985 43163
rect 26985 43129 27019 43163
rect 27019 43129 27028 43163
rect 26976 43120 27028 43129
rect 1584 43095 1636 43104
rect 1584 43061 1593 43095
rect 1593 43061 1627 43095
rect 1627 43061 1636 43095
rect 1584 43052 1636 43061
rect 2044 43052 2096 43104
rect 18236 43052 18288 43104
rect 19248 43052 19300 43104
rect 21272 43052 21324 43104
rect 27160 43052 27212 43104
rect 31944 43052 31996 43104
rect 35900 43095 35952 43104
rect 35900 43061 35909 43095
rect 35909 43061 35943 43095
rect 35943 43061 35952 43095
rect 35900 43052 35952 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 22652 42848 22704 42900
rect 20168 42780 20220 42832
rect 26240 42891 26292 42900
rect 26240 42857 26249 42891
rect 26249 42857 26283 42891
rect 26283 42857 26292 42891
rect 27068 42891 27120 42900
rect 26240 42848 26292 42857
rect 27068 42857 27077 42891
rect 27077 42857 27111 42891
rect 27111 42857 27120 42891
rect 27068 42848 27120 42857
rect 37832 42848 37884 42900
rect 1584 42712 1636 42764
rect 2780 42755 2832 42764
rect 2780 42721 2789 42755
rect 2789 42721 2823 42755
rect 2823 42721 2832 42755
rect 2780 42712 2832 42721
rect 16672 42712 16724 42764
rect 23480 42755 23532 42764
rect 23480 42721 23489 42755
rect 23489 42721 23523 42755
rect 23523 42721 23532 42755
rect 23480 42712 23532 42721
rect 23572 42712 23624 42764
rect 23940 42712 23992 42764
rect 26884 42755 26936 42764
rect 26884 42721 26893 42755
rect 26893 42721 26927 42755
rect 26927 42721 26936 42755
rect 26884 42712 26936 42721
rect 30380 42712 30432 42764
rect 30932 42712 30984 42764
rect 1584 42619 1636 42628
rect 1584 42585 1593 42619
rect 1593 42585 1627 42619
rect 1627 42585 1636 42619
rect 1584 42576 1636 42585
rect 18604 42644 18656 42696
rect 20812 42644 20864 42696
rect 21180 42687 21232 42696
rect 21180 42653 21189 42687
rect 21189 42653 21223 42687
rect 21223 42653 21232 42687
rect 21180 42644 21232 42653
rect 21456 42687 21508 42696
rect 21456 42653 21465 42687
rect 21465 42653 21499 42687
rect 21499 42653 21508 42687
rect 21456 42644 21508 42653
rect 22192 42644 22244 42696
rect 25136 42687 25188 42696
rect 25136 42653 25170 42687
rect 25170 42653 25188 42687
rect 19984 42576 20036 42628
rect 21272 42576 21324 42628
rect 25136 42644 25188 42653
rect 26976 42644 27028 42696
rect 23940 42576 23992 42628
rect 27344 42644 27396 42696
rect 29920 42644 29972 42696
rect 16488 42508 16540 42560
rect 18328 42508 18380 42560
rect 19248 42508 19300 42560
rect 20260 42551 20312 42560
rect 20260 42517 20269 42551
rect 20269 42517 20303 42551
rect 20303 42517 20312 42551
rect 20260 42508 20312 42517
rect 22284 42508 22336 42560
rect 22836 42551 22888 42560
rect 22836 42517 22845 42551
rect 22845 42517 22879 42551
rect 22879 42517 22888 42551
rect 22836 42508 22888 42517
rect 23756 42508 23808 42560
rect 29368 42576 29420 42628
rect 30012 42576 30064 42628
rect 27712 42551 27764 42560
rect 27712 42517 27721 42551
rect 27721 42517 27755 42551
rect 27755 42517 27764 42551
rect 27712 42508 27764 42517
rect 27804 42508 27856 42560
rect 29644 42508 29696 42560
rect 31944 42687 31996 42696
rect 31944 42653 31962 42687
rect 31962 42653 31996 42687
rect 31944 42644 31996 42653
rect 33048 42644 33100 42696
rect 36268 42687 36320 42696
rect 36268 42653 36277 42687
rect 36277 42653 36311 42687
rect 36311 42653 36320 42687
rect 36268 42644 36320 42653
rect 36452 42619 36504 42628
rect 36452 42585 36461 42619
rect 36461 42585 36495 42619
rect 36495 42585 36504 42619
rect 36452 42576 36504 42585
rect 38108 42619 38160 42628
rect 38108 42585 38117 42619
rect 38117 42585 38151 42619
rect 38151 42585 38160 42619
rect 38108 42576 38160 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 1584 42304 1636 42356
rect 20168 42304 20220 42356
rect 23296 42304 23348 42356
rect 24032 42304 24084 42356
rect 27804 42304 27856 42356
rect 29368 42347 29420 42356
rect 29368 42313 29377 42347
rect 29377 42313 29411 42347
rect 29411 42313 29420 42347
rect 29368 42304 29420 42313
rect 31116 42304 31168 42356
rect 36452 42304 36504 42356
rect 2044 42211 2096 42220
rect 2044 42177 2053 42211
rect 2053 42177 2087 42211
rect 2087 42177 2096 42211
rect 2044 42168 2096 42177
rect 9680 42211 9732 42220
rect 9680 42177 9689 42211
rect 9689 42177 9723 42211
rect 9723 42177 9732 42211
rect 9680 42168 9732 42177
rect 16580 42168 16632 42220
rect 18328 42211 18380 42220
rect 18328 42177 18362 42211
rect 18362 42177 18380 42211
rect 18328 42168 18380 42177
rect 20996 42211 21048 42220
rect 20996 42177 21014 42211
rect 21014 42177 21048 42211
rect 20996 42168 21048 42177
rect 27712 42236 27764 42288
rect 29920 42236 29972 42288
rect 22284 42211 22336 42220
rect 22284 42177 22293 42211
rect 22293 42177 22327 42211
rect 22327 42177 22336 42211
rect 22284 42168 22336 42177
rect 22376 42211 22428 42220
rect 22376 42177 22385 42211
rect 22385 42177 22419 42211
rect 22419 42177 22428 42211
rect 22376 42168 22428 42177
rect 22836 42168 22888 42220
rect 23756 42211 23808 42220
rect 23756 42177 23765 42211
rect 23765 42177 23799 42211
rect 23799 42177 23808 42211
rect 23756 42168 23808 42177
rect 27160 42211 27212 42220
rect 27160 42177 27169 42211
rect 27169 42177 27203 42211
rect 27203 42177 27212 42211
rect 27160 42168 27212 42177
rect 30380 42211 30432 42220
rect 2872 42100 2924 42152
rect 2964 42143 3016 42152
rect 2964 42109 2973 42143
rect 2973 42109 3007 42143
rect 3007 42109 3016 42143
rect 10416 42143 10468 42152
rect 2964 42100 3016 42109
rect 10416 42109 10425 42143
rect 10425 42109 10459 42143
rect 10459 42109 10468 42143
rect 10416 42100 10468 42109
rect 21272 42143 21324 42152
rect 21272 42109 21281 42143
rect 21281 42109 21315 42143
rect 21315 42109 21324 42143
rect 21272 42100 21324 42109
rect 22744 42143 22796 42152
rect 22744 42109 22753 42143
rect 22753 42109 22787 42143
rect 22787 42109 22796 42143
rect 22744 42100 22796 42109
rect 23296 42100 23348 42152
rect 30380 42177 30389 42211
rect 30389 42177 30423 42211
rect 30423 42177 30432 42211
rect 30380 42168 30432 42177
rect 30472 42168 30524 42220
rect 33876 42211 33928 42220
rect 33876 42177 33910 42211
rect 33910 42177 33928 42211
rect 33876 42168 33928 42177
rect 36268 42168 36320 42220
rect 37372 42168 37424 42220
rect 27712 42100 27764 42152
rect 30012 42100 30064 42152
rect 33048 42100 33100 42152
rect 14464 42032 14516 42084
rect 10416 41964 10468 42016
rect 19892 42007 19944 42016
rect 19892 41973 19901 42007
rect 19901 41973 19935 42007
rect 19935 41973 19944 42007
rect 19892 41964 19944 41973
rect 23848 42032 23900 42084
rect 22100 42007 22152 42016
rect 22100 41973 22109 42007
rect 22109 41973 22143 42007
rect 22143 41973 22152 42007
rect 22100 41964 22152 41973
rect 26976 42007 27028 42016
rect 26976 41973 26985 42007
rect 26985 41973 27019 42007
rect 27019 41973 27028 42007
rect 26976 41964 27028 41973
rect 29644 42007 29696 42016
rect 29644 41973 29653 42007
rect 29653 41973 29687 42007
rect 29687 41973 29696 42007
rect 29644 41964 29696 41973
rect 34796 41964 34848 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 2872 41803 2924 41812
rect 2872 41769 2881 41803
rect 2881 41769 2915 41803
rect 2915 41769 2924 41803
rect 2872 41760 2924 41769
rect 18604 41803 18656 41812
rect 18604 41769 18613 41803
rect 18613 41769 18647 41803
rect 18647 41769 18656 41803
rect 18604 41760 18656 41769
rect 20996 41760 21048 41812
rect 22744 41803 22796 41812
rect 22744 41769 22753 41803
rect 22753 41769 22787 41803
rect 22787 41769 22796 41803
rect 22744 41760 22796 41769
rect 33876 41760 33928 41812
rect 10048 41667 10100 41676
rect 10048 41633 10057 41667
rect 10057 41633 10091 41667
rect 10091 41633 10100 41667
rect 10048 41624 10100 41633
rect 18236 41667 18288 41676
rect 18236 41633 18245 41667
rect 18245 41633 18279 41667
rect 18279 41633 18288 41667
rect 18236 41624 18288 41633
rect 20168 41624 20220 41676
rect 23480 41624 23532 41676
rect 23848 41624 23900 41676
rect 29920 41667 29972 41676
rect 29920 41633 29929 41667
rect 29929 41633 29963 41667
rect 29963 41633 29972 41667
rect 29920 41624 29972 41633
rect 1400 41599 1452 41608
rect 1400 41565 1409 41599
rect 1409 41565 1443 41599
rect 1443 41565 1452 41599
rect 1400 41556 1452 41565
rect 8852 41556 8904 41608
rect 9680 41599 9732 41608
rect 9680 41565 9689 41599
rect 9689 41565 9723 41599
rect 9723 41565 9732 41599
rect 9680 41556 9732 41565
rect 16488 41599 16540 41608
rect 16488 41565 16522 41599
rect 16522 41565 16540 41599
rect 16488 41556 16540 41565
rect 19432 41556 19484 41608
rect 16580 41488 16632 41540
rect 8392 41420 8444 41472
rect 10048 41420 10100 41472
rect 18052 41488 18104 41540
rect 19248 41488 19300 41540
rect 23664 41556 23716 41608
rect 26976 41556 27028 41608
rect 27620 41556 27672 41608
rect 28632 41556 28684 41608
rect 30380 41556 30432 41608
rect 31208 41624 31260 41676
rect 37096 41667 37148 41676
rect 37096 41633 37105 41667
rect 37105 41633 37139 41667
rect 37139 41633 37148 41667
rect 37096 41624 37148 41633
rect 31116 41556 31168 41608
rect 34244 41556 34296 41608
rect 34520 41556 34572 41608
rect 21456 41488 21508 41540
rect 34612 41488 34664 41540
rect 37464 41488 37516 41540
rect 17592 41463 17644 41472
rect 17592 41429 17601 41463
rect 17601 41429 17635 41463
rect 17635 41429 17644 41463
rect 17592 41420 17644 41429
rect 17684 41420 17736 41472
rect 20628 41420 20680 41472
rect 26148 41420 26200 41472
rect 28908 41420 28960 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 10508 41259 10560 41268
rect 10508 41225 10517 41259
rect 10517 41225 10551 41259
rect 10551 41225 10560 41259
rect 10508 41216 10560 41225
rect 26884 41216 26936 41268
rect 27712 41216 27764 41268
rect 30012 41259 30064 41268
rect 30012 41225 30021 41259
rect 30021 41225 30055 41259
rect 30055 41225 30064 41259
rect 30012 41216 30064 41225
rect 31116 41259 31168 41268
rect 31116 41225 31125 41259
rect 31125 41225 31159 41259
rect 31159 41225 31168 41259
rect 31116 41216 31168 41225
rect 34244 41259 34296 41268
rect 9680 41148 9732 41200
rect 21272 41148 21324 41200
rect 8392 41123 8444 41132
rect 8392 41089 8401 41123
rect 8401 41089 8435 41123
rect 8435 41089 8444 41123
rect 8392 41080 8444 41089
rect 19432 41123 19484 41132
rect 19432 41089 19441 41123
rect 19441 41089 19475 41123
rect 19475 41089 19484 41123
rect 19432 41080 19484 41089
rect 21180 41080 21232 41132
rect 23388 41148 23440 41200
rect 28908 41191 28960 41200
rect 22744 41080 22796 41132
rect 20628 40876 20680 40928
rect 25228 41080 25280 41132
rect 26976 41123 27028 41132
rect 26976 41089 26985 41123
rect 26985 41089 27019 41123
rect 27019 41089 27028 41123
rect 26976 41080 27028 41089
rect 28908 41157 28942 41191
rect 28942 41157 28960 41191
rect 28908 41148 28960 41157
rect 30932 41123 30984 41132
rect 30932 41089 30941 41123
rect 30941 41089 30975 41123
rect 30975 41089 30984 41123
rect 30932 41080 30984 41089
rect 24860 40944 24912 40996
rect 27988 41012 28040 41064
rect 28632 41055 28684 41064
rect 28632 41021 28641 41055
rect 28641 41021 28675 41055
rect 28675 41021 28684 41055
rect 28632 41012 28684 41021
rect 31760 41012 31812 41064
rect 33048 41148 33100 41200
rect 34244 41225 34253 41259
rect 34253 41225 34287 41259
rect 34287 41225 34296 41259
rect 34244 41216 34296 41225
rect 37464 41259 37516 41268
rect 37464 41225 37473 41259
rect 37473 41225 37507 41259
rect 37507 41225 37516 41259
rect 37464 41216 37516 41225
rect 32680 41123 32732 41132
rect 32680 41089 32714 41123
rect 32714 41089 32732 41123
rect 32680 41080 32732 41089
rect 35992 41080 36044 41132
rect 34796 41012 34848 41064
rect 35348 41012 35400 41064
rect 25136 40876 25188 40928
rect 26884 40876 26936 40928
rect 38384 40944 38436 40996
rect 35808 40876 35860 40928
rect 36084 40919 36136 40928
rect 36084 40885 36093 40919
rect 36093 40885 36127 40919
rect 36127 40885 36136 40919
rect 36084 40876 36136 40885
rect 36268 40876 36320 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 21272 40672 21324 40724
rect 23664 40672 23716 40724
rect 26056 40672 26108 40724
rect 32680 40715 32732 40724
rect 32680 40681 32689 40715
rect 32689 40681 32723 40715
rect 32723 40681 32732 40715
rect 32680 40672 32732 40681
rect 34520 40672 34572 40724
rect 34704 40672 34756 40724
rect 10968 40536 11020 40588
rect 15292 40536 15344 40588
rect 18696 40536 18748 40588
rect 24860 40536 24912 40588
rect 25872 40604 25924 40656
rect 26148 40604 26200 40656
rect 34612 40536 34664 40588
rect 36268 40579 36320 40588
rect 36268 40545 36277 40579
rect 36277 40545 36311 40579
rect 36311 40545 36320 40579
rect 36268 40536 36320 40545
rect 38200 40536 38252 40588
rect 1584 40511 1636 40520
rect 1584 40477 1593 40511
rect 1593 40477 1627 40511
rect 1627 40477 1636 40511
rect 1584 40468 1636 40477
rect 9680 40511 9732 40520
rect 9680 40477 9689 40511
rect 9689 40477 9723 40511
rect 9723 40477 9732 40511
rect 9680 40468 9732 40477
rect 16764 40468 16816 40520
rect 21180 40468 21232 40520
rect 23664 40511 23716 40520
rect 23664 40477 23673 40511
rect 23673 40477 23707 40511
rect 23707 40477 23716 40511
rect 23664 40468 23716 40477
rect 21088 40443 21140 40452
rect 21088 40409 21097 40443
rect 21097 40409 21131 40443
rect 21131 40409 21140 40443
rect 21088 40400 21140 40409
rect 22100 40400 22152 40452
rect 16672 40375 16724 40384
rect 16672 40341 16681 40375
rect 16681 40341 16715 40375
rect 16715 40341 16724 40375
rect 16672 40332 16724 40341
rect 27712 40511 27764 40520
rect 27712 40477 27730 40511
rect 27730 40477 27764 40511
rect 27988 40511 28040 40520
rect 27712 40468 27764 40477
rect 27988 40477 27997 40511
rect 27997 40477 28031 40511
rect 28031 40477 28040 40511
rect 27988 40468 28040 40477
rect 32864 40511 32916 40520
rect 32864 40477 32873 40511
rect 32873 40477 32907 40511
rect 32907 40477 32916 40511
rect 32864 40468 32916 40477
rect 34796 40468 34848 40520
rect 35808 40511 35860 40520
rect 35808 40477 35817 40511
rect 35817 40477 35851 40511
rect 35851 40477 35860 40511
rect 35808 40468 35860 40477
rect 24952 40400 25004 40452
rect 25228 40400 25280 40452
rect 35348 40400 35400 40452
rect 37372 40400 37424 40452
rect 25596 40375 25648 40384
rect 25596 40341 25605 40375
rect 25605 40341 25639 40375
rect 25639 40341 25648 40375
rect 25596 40332 25648 40341
rect 25780 40332 25832 40384
rect 33600 40332 33652 40384
rect 35624 40375 35676 40384
rect 35624 40341 35633 40375
rect 35633 40341 35667 40375
rect 35667 40341 35676 40375
rect 35624 40332 35676 40341
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 9772 40128 9824 40180
rect 3424 40103 3476 40112
rect 3424 40069 3433 40103
rect 3433 40069 3467 40103
rect 3467 40069 3476 40103
rect 3424 40060 3476 40069
rect 9680 40060 9732 40112
rect 1584 40035 1636 40044
rect 1584 40001 1593 40035
rect 1593 40001 1627 40035
rect 1627 40001 1636 40035
rect 1584 39992 1636 40001
rect 16672 40060 16724 40112
rect 17868 40128 17920 40180
rect 20352 40128 20404 40180
rect 23664 40128 23716 40180
rect 22652 40060 22704 40112
rect 26976 40128 27028 40180
rect 30656 40128 30708 40180
rect 30748 40103 30800 40112
rect 18144 39992 18196 40044
rect 20352 40035 20404 40044
rect 20352 40001 20361 40035
rect 20361 40001 20395 40035
rect 20395 40001 20404 40035
rect 20352 39992 20404 40001
rect 1768 39967 1820 39976
rect 1768 39933 1777 39967
rect 1777 39933 1811 39967
rect 1811 39933 1820 39967
rect 1768 39924 1820 39933
rect 19524 39924 19576 39976
rect 21180 39992 21232 40044
rect 21916 39992 21968 40044
rect 24860 39992 24912 40044
rect 25780 40035 25832 40044
rect 25780 40001 25789 40035
rect 25789 40001 25823 40035
rect 25823 40001 25832 40035
rect 25780 39992 25832 40001
rect 25872 39992 25924 40044
rect 30748 40069 30757 40103
rect 30757 40069 30791 40103
rect 30791 40069 30800 40103
rect 30748 40060 30800 40069
rect 27988 39992 28040 40044
rect 20628 39924 20680 39976
rect 20996 39924 21048 39976
rect 23664 39924 23716 39976
rect 21272 39856 21324 39908
rect 24952 39856 25004 39908
rect 20812 39788 20864 39840
rect 24676 39831 24728 39840
rect 24676 39797 24685 39831
rect 24685 39797 24719 39831
rect 24719 39797 24728 39831
rect 24676 39788 24728 39797
rect 25780 39831 25832 39840
rect 25780 39797 25789 39831
rect 25789 39797 25823 39831
rect 25823 39797 25832 39831
rect 25780 39788 25832 39797
rect 28908 39992 28960 40044
rect 31576 40035 31628 40044
rect 31576 40001 31585 40035
rect 31585 40001 31619 40035
rect 31619 40001 31628 40035
rect 31576 39992 31628 40001
rect 31760 39992 31812 40044
rect 33232 40035 33284 40044
rect 33232 40001 33250 40035
rect 33250 40001 33284 40035
rect 33232 39992 33284 40001
rect 34244 40035 34296 40044
rect 34244 40001 34278 40035
rect 34278 40001 34296 40035
rect 34244 39992 34296 40001
rect 34704 39992 34756 40044
rect 35992 40035 36044 40044
rect 33968 39967 34020 39976
rect 33968 39933 33977 39967
rect 33977 39933 34011 39967
rect 34011 39933 34020 39967
rect 33968 39924 34020 39933
rect 35992 40001 36001 40035
rect 36001 40001 36035 40035
rect 36035 40001 36044 40035
rect 35992 39992 36044 40001
rect 37372 40035 37424 40044
rect 37372 40001 37381 40035
rect 37381 40001 37415 40035
rect 37415 40001 37424 40035
rect 37372 39992 37424 40001
rect 37924 39924 37976 39976
rect 31392 39831 31444 39840
rect 31392 39797 31401 39831
rect 31401 39797 31435 39831
rect 31435 39797 31444 39831
rect 31392 39788 31444 39797
rect 32128 39831 32180 39840
rect 32128 39797 32137 39831
rect 32137 39797 32171 39831
rect 32171 39797 32180 39831
rect 32128 39788 32180 39797
rect 35348 39831 35400 39840
rect 35348 39797 35357 39831
rect 35357 39797 35391 39831
rect 35391 39797 35400 39831
rect 35348 39788 35400 39797
rect 35808 39831 35860 39840
rect 35808 39797 35817 39831
rect 35817 39797 35851 39831
rect 35851 39797 35860 39831
rect 35808 39788 35860 39797
rect 38200 39788 38252 39840
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 1768 39584 1820 39636
rect 16764 39627 16816 39636
rect 16764 39593 16773 39627
rect 16773 39593 16807 39627
rect 16807 39593 16816 39627
rect 16764 39584 16816 39593
rect 18144 39627 18196 39636
rect 18144 39593 18153 39627
rect 18153 39593 18187 39627
rect 18187 39593 18196 39627
rect 18144 39584 18196 39593
rect 25044 39584 25096 39636
rect 25596 39584 25648 39636
rect 28908 39584 28960 39636
rect 31576 39584 31628 39636
rect 32864 39584 32916 39636
rect 33232 39584 33284 39636
rect 34244 39584 34296 39636
rect 17592 39448 17644 39500
rect 21272 39448 21324 39500
rect 2136 39423 2188 39432
rect 2136 39389 2145 39423
rect 2145 39389 2179 39423
rect 2179 39389 2188 39423
rect 2136 39380 2188 39389
rect 16856 39312 16908 39364
rect 18328 39380 18380 39432
rect 18696 39312 18748 39364
rect 20904 39355 20956 39364
rect 20904 39321 20922 39355
rect 20922 39321 20956 39355
rect 20904 39312 20956 39321
rect 21916 39423 21968 39432
rect 21916 39389 21925 39423
rect 21925 39389 21959 39423
rect 21959 39389 21968 39423
rect 21916 39380 21968 39389
rect 24676 39380 24728 39432
rect 25780 39448 25832 39500
rect 30656 39448 30708 39500
rect 25136 39423 25188 39432
rect 25136 39389 25145 39423
rect 25145 39389 25179 39423
rect 25179 39389 25188 39423
rect 28356 39423 28408 39432
rect 25136 39380 25188 39389
rect 28356 39389 28365 39423
rect 28365 39389 28399 39423
rect 28399 39389 28408 39423
rect 28356 39380 28408 39389
rect 32128 39423 32180 39432
rect 29552 39312 29604 39364
rect 32128 39389 32137 39423
rect 32137 39389 32171 39423
rect 32171 39389 32180 39423
rect 32128 39380 32180 39389
rect 32312 39380 32364 39432
rect 32496 39380 32548 39432
rect 35808 39584 35860 39636
rect 34796 39516 34848 39568
rect 34704 39448 34756 39500
rect 36084 39448 36136 39500
rect 38108 39491 38160 39500
rect 38108 39457 38117 39491
rect 38117 39457 38151 39491
rect 38151 39457 38160 39491
rect 38108 39448 38160 39457
rect 34612 39312 34664 39364
rect 20076 39244 20128 39296
rect 21824 39244 21876 39296
rect 25320 39287 25372 39296
rect 25320 39253 25329 39287
rect 25329 39253 25363 39287
rect 25363 39253 25372 39287
rect 25320 39244 25372 39253
rect 34704 39287 34756 39296
rect 34704 39253 34713 39287
rect 34713 39253 34747 39287
rect 34747 39253 34756 39287
rect 34704 39244 34756 39253
rect 36452 39355 36504 39364
rect 34980 39287 35032 39296
rect 34980 39253 34989 39287
rect 34989 39253 35023 39287
rect 35023 39253 35032 39287
rect 34980 39244 35032 39253
rect 36452 39321 36461 39355
rect 36461 39321 36495 39355
rect 36495 39321 36504 39355
rect 36452 39312 36504 39321
rect 35348 39244 35400 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 18328 39083 18380 39092
rect 18328 39049 18337 39083
rect 18337 39049 18371 39083
rect 18371 39049 18380 39083
rect 18328 39040 18380 39049
rect 20904 39040 20956 39092
rect 28356 39040 28408 39092
rect 32496 39083 32548 39092
rect 32496 39049 32505 39083
rect 32505 39049 32539 39083
rect 32539 39049 32548 39083
rect 32496 39040 32548 39049
rect 36452 39040 36504 39092
rect 1676 38972 1728 39024
rect 16856 38947 16908 38956
rect 16856 38913 16865 38947
rect 16865 38913 16899 38947
rect 16899 38913 16908 38947
rect 16856 38904 16908 38913
rect 19432 38972 19484 39024
rect 18604 38947 18656 38956
rect 18604 38913 18613 38947
rect 18613 38913 18647 38947
rect 18647 38913 18656 38947
rect 19984 38947 20036 38956
rect 18604 38904 18656 38913
rect 19984 38913 19993 38947
rect 19993 38913 20027 38947
rect 20027 38913 20036 38947
rect 19984 38904 20036 38913
rect 20168 38947 20220 38956
rect 20168 38913 20177 38947
rect 20177 38913 20211 38947
rect 20211 38913 20220 38947
rect 20168 38904 20220 38913
rect 20812 38947 20864 38956
rect 20812 38913 20821 38947
rect 20821 38913 20855 38947
rect 20855 38913 20864 38947
rect 20812 38904 20864 38913
rect 21732 38904 21784 38956
rect 24676 38904 24728 38956
rect 25044 38947 25096 38956
rect 25044 38913 25053 38947
rect 25053 38913 25087 38947
rect 25087 38913 25096 38947
rect 25044 38904 25096 38913
rect 1860 38879 1912 38888
rect 1860 38845 1869 38879
rect 1869 38845 1903 38879
rect 1903 38845 1912 38879
rect 1860 38836 1912 38845
rect 2780 38836 2832 38888
rect 2872 38879 2924 38888
rect 2872 38845 2881 38879
rect 2881 38845 2915 38879
rect 2915 38845 2924 38879
rect 2872 38836 2924 38845
rect 17868 38836 17920 38888
rect 21824 38879 21876 38888
rect 21824 38845 21833 38879
rect 21833 38845 21867 38879
rect 21867 38845 21876 38879
rect 21824 38836 21876 38845
rect 25412 38904 25464 38956
rect 25780 38947 25832 38956
rect 25780 38913 25789 38947
rect 25789 38913 25823 38947
rect 25823 38913 25832 38947
rect 25780 38904 25832 38913
rect 26056 38947 26108 38956
rect 26056 38913 26065 38947
rect 26065 38913 26099 38947
rect 26099 38913 26108 38947
rect 26056 38904 26108 38913
rect 31760 38972 31812 39024
rect 35624 39015 35676 39024
rect 35624 38981 35658 39015
rect 35658 38981 35676 39015
rect 35624 38972 35676 38981
rect 31392 38904 31444 38956
rect 31852 38904 31904 38956
rect 32312 38947 32364 38956
rect 32312 38913 32321 38947
rect 32321 38913 32355 38947
rect 32355 38913 32364 38947
rect 32312 38904 32364 38913
rect 33968 38904 34020 38956
rect 37464 38947 37516 38956
rect 37464 38913 37473 38947
rect 37473 38913 37507 38947
rect 37507 38913 37516 38947
rect 37464 38904 37516 38913
rect 25228 38836 25280 38888
rect 32128 38879 32180 38888
rect 32128 38845 32137 38879
rect 32137 38845 32171 38879
rect 32171 38845 32180 38879
rect 32128 38836 32180 38845
rect 25136 38768 25188 38820
rect 34980 38768 35032 38820
rect 14096 38743 14148 38752
rect 14096 38709 14105 38743
rect 14105 38709 14139 38743
rect 14139 38709 14148 38743
rect 14096 38700 14148 38709
rect 16580 38700 16632 38752
rect 20904 38700 20956 38752
rect 23940 38700 23992 38752
rect 25872 38700 25924 38752
rect 32312 38700 32364 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 1860 38539 1912 38548
rect 1860 38505 1869 38539
rect 1869 38505 1903 38539
rect 1903 38505 1912 38539
rect 1860 38496 1912 38505
rect 2780 38539 2832 38548
rect 2780 38505 2789 38539
rect 2789 38505 2823 38539
rect 2823 38505 2832 38539
rect 2780 38496 2832 38505
rect 17592 38539 17644 38548
rect 17592 38505 17601 38539
rect 17601 38505 17635 38539
rect 17635 38505 17644 38539
rect 17592 38496 17644 38505
rect 19984 38496 20036 38548
rect 20352 38539 20404 38548
rect 20352 38505 20361 38539
rect 20361 38505 20395 38539
rect 20395 38505 20404 38539
rect 20352 38496 20404 38505
rect 32312 38539 32364 38548
rect 32312 38505 32321 38539
rect 32321 38505 32355 38539
rect 32355 38505 32364 38539
rect 32312 38496 32364 38505
rect 20168 38428 20220 38480
rect 24860 38428 24912 38480
rect 26056 38428 26108 38480
rect 18144 38360 18196 38412
rect 18604 38360 18656 38412
rect 20352 38360 20404 38412
rect 20628 38360 20680 38412
rect 4712 38292 4764 38344
rect 16488 38292 16540 38344
rect 17868 38335 17920 38344
rect 17868 38301 17877 38335
rect 17877 38301 17911 38335
rect 17911 38301 17920 38335
rect 17868 38292 17920 38301
rect 20076 38335 20128 38344
rect 20076 38301 20085 38335
rect 20085 38301 20119 38335
rect 20119 38301 20128 38335
rect 21272 38360 21324 38412
rect 25228 38360 25280 38412
rect 32128 38360 32180 38412
rect 37096 38403 37148 38412
rect 37096 38369 37105 38403
rect 37105 38369 37139 38403
rect 37139 38369 37148 38403
rect 37096 38360 37148 38369
rect 38200 38360 38252 38412
rect 20076 38292 20128 38301
rect 24676 38335 24728 38344
rect 24676 38301 24685 38335
rect 24685 38301 24719 38335
rect 24719 38301 24728 38335
rect 24860 38335 24912 38344
rect 24676 38292 24728 38301
rect 24860 38301 24869 38335
rect 24869 38301 24903 38335
rect 24903 38301 24912 38335
rect 24860 38292 24912 38301
rect 15936 38224 15988 38276
rect 17500 38156 17552 38208
rect 20444 38224 20496 38276
rect 23020 38224 23072 38276
rect 27988 38292 28040 38344
rect 30656 38292 30708 38344
rect 31668 38292 31720 38344
rect 33600 38335 33652 38344
rect 33600 38301 33609 38335
rect 33609 38301 33643 38335
rect 33643 38301 33652 38335
rect 33600 38292 33652 38301
rect 35440 38335 35492 38344
rect 35440 38301 35449 38335
rect 35449 38301 35483 38335
rect 35483 38301 35492 38335
rect 35440 38292 35492 38301
rect 35900 38292 35952 38344
rect 21180 38199 21232 38208
rect 21180 38165 21189 38199
rect 21189 38165 21223 38199
rect 21223 38165 21232 38199
rect 21180 38156 21232 38165
rect 27712 38267 27764 38276
rect 27712 38233 27746 38267
rect 27746 38233 27764 38267
rect 27712 38224 27764 38233
rect 32220 38224 32272 38276
rect 24216 38156 24268 38208
rect 24860 38156 24912 38208
rect 27528 38156 27580 38208
rect 37464 38224 37516 38276
rect 33140 38156 33192 38208
rect 35808 38199 35860 38208
rect 35808 38165 35817 38199
rect 35817 38165 35851 38199
rect 35851 38165 35860 38199
rect 35808 38156 35860 38165
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 15936 37995 15988 38004
rect 15936 37961 15945 37995
rect 15945 37961 15979 37995
rect 15979 37961 15988 37995
rect 15936 37952 15988 37961
rect 17776 37952 17828 38004
rect 18144 37952 18196 38004
rect 20260 37995 20312 38004
rect 20260 37961 20269 37995
rect 20269 37961 20303 37995
rect 20303 37961 20312 37995
rect 20260 37952 20312 37961
rect 27712 37952 27764 38004
rect 29828 37995 29880 38004
rect 17500 37884 17552 37936
rect 20444 37927 20496 37936
rect 14096 37859 14148 37868
rect 14096 37825 14105 37859
rect 14105 37825 14139 37859
rect 14139 37825 14148 37859
rect 14096 37816 14148 37825
rect 16580 37816 16632 37868
rect 16764 37816 16816 37868
rect 18696 37859 18748 37868
rect 18696 37825 18705 37859
rect 18705 37825 18739 37859
rect 18739 37825 18748 37859
rect 18696 37816 18748 37825
rect 20444 37893 20453 37927
rect 20453 37893 20487 37927
rect 20487 37893 20496 37927
rect 20444 37884 20496 37893
rect 24860 37927 24912 37936
rect 24860 37893 24869 37927
rect 24869 37893 24903 37927
rect 24903 37893 24912 37927
rect 24860 37884 24912 37893
rect 25320 37884 25372 37936
rect 27528 37884 27580 37936
rect 19524 37859 19576 37868
rect 19524 37825 19533 37859
rect 19533 37825 19567 37859
rect 19567 37825 19576 37859
rect 19524 37816 19576 37825
rect 20076 37859 20128 37868
rect 20076 37825 20085 37859
rect 20085 37825 20119 37859
rect 20119 37825 20128 37859
rect 20076 37816 20128 37825
rect 20352 37859 20404 37868
rect 20352 37825 20361 37859
rect 20361 37825 20395 37859
rect 20395 37825 20404 37859
rect 20352 37816 20404 37825
rect 21180 37816 21232 37868
rect 23112 37859 23164 37868
rect 23112 37825 23121 37859
rect 23121 37825 23155 37859
rect 23155 37825 23164 37859
rect 23112 37816 23164 37825
rect 23940 37859 23992 37868
rect 23940 37825 23949 37859
rect 23949 37825 23983 37859
rect 23983 37825 23992 37859
rect 23940 37816 23992 37825
rect 24124 37859 24176 37868
rect 24124 37825 24133 37859
rect 24133 37825 24167 37859
rect 24167 37825 24176 37859
rect 24124 37816 24176 37825
rect 24216 37859 24268 37868
rect 24216 37825 24225 37859
rect 24225 37825 24259 37859
rect 24259 37825 24268 37859
rect 24216 37816 24268 37825
rect 26792 37816 26844 37868
rect 16488 37748 16540 37800
rect 27344 37859 27396 37868
rect 27344 37825 27353 37859
rect 27353 37825 27387 37859
rect 27387 37825 27396 37859
rect 28908 37859 28960 37868
rect 27344 37816 27396 37825
rect 28908 37825 28917 37859
rect 28917 37825 28951 37859
rect 28951 37825 28960 37859
rect 28908 37816 28960 37825
rect 29828 37961 29837 37995
rect 29837 37961 29871 37995
rect 29871 37961 29880 37995
rect 29828 37952 29880 37961
rect 32312 37952 32364 38004
rect 37464 37995 37516 38004
rect 37464 37961 37473 37995
rect 37473 37961 37507 37995
rect 37507 37961 37516 37995
rect 37464 37952 37516 37961
rect 32128 37884 32180 37936
rect 30104 37816 30156 37868
rect 32220 37816 32272 37868
rect 34520 37859 34572 37868
rect 34520 37825 34529 37859
rect 34529 37825 34563 37859
rect 34563 37825 34572 37859
rect 34520 37816 34572 37825
rect 35624 37859 35676 37868
rect 35624 37825 35658 37859
rect 35658 37825 35676 37859
rect 35624 37816 35676 37825
rect 37280 37816 37332 37868
rect 38292 37816 38344 37868
rect 29000 37791 29052 37800
rect 29000 37757 29009 37791
rect 29009 37757 29043 37791
rect 29043 37757 29052 37791
rect 29000 37748 29052 37757
rect 31668 37748 31720 37800
rect 35348 37791 35400 37800
rect 35348 37757 35357 37791
rect 35357 37757 35391 37791
rect 35391 37757 35400 37791
rect 35348 37748 35400 37757
rect 27252 37680 27304 37732
rect 14648 37612 14700 37664
rect 18512 37655 18564 37664
rect 18512 37621 18521 37655
rect 18521 37621 18555 37655
rect 18555 37621 18564 37655
rect 18512 37612 18564 37621
rect 19340 37655 19392 37664
rect 19340 37621 19349 37655
rect 19349 37621 19383 37655
rect 19383 37621 19392 37655
rect 19340 37612 19392 37621
rect 20720 37612 20772 37664
rect 21272 37655 21324 37664
rect 21272 37621 21281 37655
rect 21281 37621 21315 37655
rect 21315 37621 21324 37655
rect 21272 37612 21324 37621
rect 23572 37612 23624 37664
rect 23664 37612 23716 37664
rect 24768 37655 24820 37664
rect 24768 37621 24777 37655
rect 24777 37621 24811 37655
rect 24811 37621 24820 37655
rect 24768 37612 24820 37621
rect 25412 37612 25464 37664
rect 30012 37655 30064 37664
rect 30012 37621 30021 37655
rect 30021 37621 30055 37655
rect 30055 37621 30064 37655
rect 30012 37612 30064 37621
rect 32772 37612 32824 37664
rect 34336 37655 34388 37664
rect 34336 37621 34345 37655
rect 34345 37621 34379 37655
rect 34379 37621 34388 37655
rect 34336 37612 34388 37621
rect 36728 37655 36780 37664
rect 36728 37621 36737 37655
rect 36737 37621 36771 37655
rect 36771 37621 36780 37655
rect 36728 37612 36780 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 16764 37451 16816 37460
rect 16764 37417 16773 37451
rect 16773 37417 16807 37451
rect 16807 37417 16816 37451
rect 16764 37408 16816 37417
rect 23020 37451 23072 37460
rect 23020 37417 23029 37451
rect 23029 37417 23063 37451
rect 23063 37417 23072 37451
rect 23020 37408 23072 37417
rect 23112 37408 23164 37460
rect 27252 37451 27304 37460
rect 27252 37417 27261 37451
rect 27261 37417 27295 37451
rect 27295 37417 27304 37451
rect 27252 37408 27304 37417
rect 29000 37451 29052 37460
rect 29000 37417 29009 37451
rect 29009 37417 29043 37451
rect 29043 37417 29052 37451
rect 29000 37408 29052 37417
rect 34520 37408 34572 37460
rect 35624 37451 35676 37460
rect 35624 37417 35633 37451
rect 35633 37417 35667 37451
rect 35667 37417 35676 37451
rect 35624 37408 35676 37417
rect 4712 37340 4764 37392
rect 10968 37340 11020 37392
rect 17868 37340 17920 37392
rect 3332 37272 3384 37324
rect 14280 37272 14332 37324
rect 20628 37272 20680 37324
rect 16488 37204 16540 37256
rect 18512 37204 18564 37256
rect 19432 37247 19484 37256
rect 19432 37213 19441 37247
rect 19441 37213 19475 37247
rect 19475 37213 19484 37247
rect 19432 37204 19484 37213
rect 14648 37179 14700 37188
rect 14648 37145 14682 37179
rect 14682 37145 14700 37179
rect 14648 37136 14700 37145
rect 17592 37136 17644 37188
rect 17776 37179 17828 37188
rect 17776 37145 17785 37179
rect 17785 37145 17819 37179
rect 17819 37145 17828 37179
rect 17776 37136 17828 37145
rect 19524 37136 19576 37188
rect 16856 37068 16908 37120
rect 17500 37068 17552 37120
rect 20260 37204 20312 37256
rect 22376 37247 22428 37256
rect 22376 37213 22385 37247
rect 22385 37213 22419 37247
rect 22419 37213 22428 37247
rect 22376 37204 22428 37213
rect 22468 37204 22520 37256
rect 22836 37272 22888 37324
rect 23572 37204 23624 37256
rect 24768 37272 24820 37324
rect 25228 37272 25280 37324
rect 27528 37340 27580 37392
rect 21272 37136 21324 37188
rect 23756 37136 23808 37188
rect 24124 37136 24176 37188
rect 25320 37204 25372 37256
rect 26240 37247 26292 37256
rect 25688 37136 25740 37188
rect 26240 37213 26249 37247
rect 26249 37213 26283 37247
rect 26283 37213 26292 37247
rect 26240 37204 26292 37213
rect 27068 37272 27120 37324
rect 27160 37204 27212 37256
rect 27712 37247 27764 37256
rect 27712 37213 27721 37247
rect 27721 37213 27755 37247
rect 27755 37213 27764 37247
rect 27712 37204 27764 37213
rect 32312 37272 32364 37324
rect 33232 37315 33284 37324
rect 33232 37281 33241 37315
rect 33241 37281 33275 37315
rect 33275 37281 33284 37315
rect 33232 37272 33284 37281
rect 36728 37272 36780 37324
rect 38108 37315 38160 37324
rect 38108 37281 38117 37315
rect 38117 37281 38151 37315
rect 38151 37281 38160 37315
rect 38108 37272 38160 37281
rect 20444 37068 20496 37120
rect 23480 37111 23532 37120
rect 23480 37077 23489 37111
rect 23489 37077 23523 37111
rect 23523 37077 23532 37111
rect 23480 37068 23532 37077
rect 25320 37111 25372 37120
rect 25320 37077 25329 37111
rect 25329 37077 25363 37111
rect 25363 37077 25372 37111
rect 25320 37068 25372 37077
rect 31760 37204 31812 37256
rect 31852 37247 31904 37256
rect 31852 37213 31861 37247
rect 31861 37213 31895 37247
rect 31895 37213 31904 37247
rect 32772 37247 32824 37256
rect 31852 37204 31904 37213
rect 32772 37213 32781 37247
rect 32781 37213 32815 37247
rect 32815 37213 32824 37247
rect 32772 37204 32824 37213
rect 33140 37204 33192 37256
rect 34520 37204 34572 37256
rect 35808 37247 35860 37256
rect 30012 37136 30064 37188
rect 30840 37068 30892 37120
rect 31392 37068 31444 37120
rect 32588 37111 32640 37120
rect 32588 37077 32597 37111
rect 32597 37077 32631 37111
rect 32631 37077 32640 37111
rect 32588 37068 32640 37077
rect 32956 37179 33008 37188
rect 32956 37145 32965 37179
rect 32965 37145 32999 37179
rect 32999 37145 33008 37179
rect 35808 37213 35817 37247
rect 35817 37213 35851 37247
rect 35851 37213 35860 37247
rect 35808 37204 35860 37213
rect 36268 37247 36320 37256
rect 36268 37213 36277 37247
rect 36277 37213 36311 37247
rect 36311 37213 36320 37247
rect 36268 37204 36320 37213
rect 32956 37136 33008 37145
rect 35992 37136 36044 37188
rect 37464 37136 37516 37188
rect 34704 37068 34756 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 20352 36864 20404 36916
rect 22468 36864 22520 36916
rect 23480 36864 23532 36916
rect 27160 36907 27212 36916
rect 27160 36873 27169 36907
rect 27169 36873 27203 36907
rect 27203 36873 27212 36907
rect 27160 36864 27212 36873
rect 28908 36864 28960 36916
rect 30104 36864 30156 36916
rect 32128 36907 32180 36916
rect 32128 36873 32137 36907
rect 32137 36873 32171 36907
rect 32171 36873 32180 36907
rect 32128 36864 32180 36873
rect 32772 36864 32824 36916
rect 35440 36864 35492 36916
rect 37464 36907 37516 36916
rect 37464 36873 37473 36907
rect 37473 36873 37507 36907
rect 37507 36873 37516 36907
rect 37464 36864 37516 36873
rect 14280 36839 14332 36848
rect 14280 36805 14289 36839
rect 14289 36805 14323 36839
rect 14323 36805 14332 36839
rect 14280 36796 14332 36805
rect 16488 36728 16540 36780
rect 20260 36796 20312 36848
rect 20720 36839 20772 36848
rect 20720 36805 20729 36839
rect 20729 36805 20763 36839
rect 20763 36805 20772 36839
rect 20720 36796 20772 36805
rect 20904 36839 20956 36848
rect 20904 36805 20939 36839
rect 20939 36805 20956 36839
rect 20904 36796 20956 36805
rect 19340 36728 19392 36780
rect 20628 36771 20680 36780
rect 20628 36737 20637 36771
rect 20637 36737 20671 36771
rect 20671 36737 20680 36771
rect 20628 36728 20680 36737
rect 23388 36796 23440 36848
rect 25412 36796 25464 36848
rect 26240 36796 26292 36848
rect 26976 36796 27028 36848
rect 23572 36771 23624 36780
rect 14372 36660 14424 36712
rect 15752 36592 15804 36644
rect 20720 36660 20772 36712
rect 23572 36737 23581 36771
rect 23581 36737 23615 36771
rect 23615 36737 23624 36771
rect 23572 36728 23624 36737
rect 23756 36771 23808 36780
rect 23756 36737 23765 36771
rect 23765 36737 23799 36771
rect 23799 36737 23808 36771
rect 23756 36728 23808 36737
rect 24952 36728 25004 36780
rect 25320 36771 25372 36780
rect 25320 36737 25329 36771
rect 25329 36737 25363 36771
rect 25363 36737 25372 36771
rect 25320 36728 25372 36737
rect 27068 36771 27120 36780
rect 27068 36737 27077 36771
rect 27077 36737 27111 36771
rect 27111 36737 27120 36771
rect 27068 36728 27120 36737
rect 30748 36796 30800 36848
rect 31760 36796 31812 36848
rect 32864 36796 32916 36848
rect 34336 36796 34388 36848
rect 30840 36728 30892 36780
rect 31576 36728 31628 36780
rect 36268 36728 36320 36780
rect 37372 36771 37424 36780
rect 37372 36737 37381 36771
rect 37381 36737 37415 36771
rect 37415 36737 37424 36771
rect 37372 36728 37424 36737
rect 38476 36728 38528 36780
rect 29552 36660 29604 36712
rect 30196 36660 30248 36712
rect 20904 36592 20956 36644
rect 26056 36592 26108 36644
rect 29644 36592 29696 36644
rect 20444 36567 20496 36576
rect 20444 36533 20453 36567
rect 20453 36533 20487 36567
rect 20487 36533 20496 36567
rect 20444 36524 20496 36533
rect 23388 36524 23440 36576
rect 26608 36524 26660 36576
rect 27344 36524 27396 36576
rect 30196 36524 30248 36576
rect 32772 36524 32824 36576
rect 32864 36524 32916 36576
rect 34612 36524 34664 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 14372 36363 14424 36372
rect 14372 36329 14381 36363
rect 14381 36329 14415 36363
rect 14415 36329 14424 36363
rect 14372 36320 14424 36329
rect 20260 36363 20312 36372
rect 20260 36329 20269 36363
rect 20269 36329 20303 36363
rect 20303 36329 20312 36363
rect 20260 36320 20312 36329
rect 19248 36252 19300 36304
rect 37372 36320 37424 36372
rect 21640 36252 21692 36304
rect 22376 36252 22428 36304
rect 24676 36295 24728 36304
rect 24676 36261 24685 36295
rect 24685 36261 24719 36295
rect 24719 36261 24728 36295
rect 24676 36252 24728 36261
rect 26976 36295 27028 36304
rect 26976 36261 26985 36295
rect 26985 36261 27019 36295
rect 27019 36261 27028 36295
rect 26976 36252 27028 36261
rect 31576 36295 31628 36304
rect 31576 36261 31585 36295
rect 31585 36261 31619 36295
rect 31619 36261 31628 36295
rect 31576 36252 31628 36261
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 3240 36159 3292 36168
rect 3240 36125 3249 36159
rect 3249 36125 3283 36159
rect 3283 36125 3292 36159
rect 3240 36116 3292 36125
rect 14096 36116 14148 36168
rect 21088 36184 21140 36236
rect 26240 36184 26292 36236
rect 21824 36116 21876 36168
rect 23848 36116 23900 36168
rect 24400 36159 24452 36168
rect 24400 36125 24409 36159
rect 24409 36125 24443 36159
rect 24443 36125 24452 36159
rect 24400 36116 24452 36125
rect 25872 36159 25924 36168
rect 25872 36125 25881 36159
rect 25881 36125 25915 36159
rect 25915 36125 25924 36159
rect 25872 36116 25924 36125
rect 27160 36159 27212 36168
rect 27160 36125 27169 36159
rect 27169 36125 27203 36159
rect 27203 36125 27212 36159
rect 27160 36116 27212 36125
rect 27528 36116 27580 36168
rect 29276 36116 29328 36168
rect 31392 36159 31444 36168
rect 31392 36125 31401 36159
rect 31401 36125 31435 36159
rect 31435 36125 31444 36159
rect 31392 36116 31444 36125
rect 35348 36116 35400 36168
rect 36176 36116 36228 36168
rect 3056 36091 3108 36100
rect 3056 36057 3065 36091
rect 3065 36057 3099 36091
rect 3099 36057 3108 36091
rect 3056 36048 3108 36057
rect 24584 36048 24636 36100
rect 36360 36048 36412 36100
rect 20720 35980 20772 36032
rect 24308 35980 24360 36032
rect 24860 35980 24912 36032
rect 37464 35980 37516 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 3056 35776 3108 35828
rect 24032 35776 24084 35828
rect 20444 35708 20496 35760
rect 23664 35708 23716 35760
rect 24492 35708 24544 35760
rect 14096 35640 14148 35692
rect 17408 35683 17460 35692
rect 17408 35649 17417 35683
rect 17417 35649 17451 35683
rect 17451 35649 17460 35683
rect 17408 35640 17460 35649
rect 23112 35683 23164 35692
rect 23112 35649 23121 35683
rect 23121 35649 23155 35683
rect 23155 35649 23164 35683
rect 23112 35640 23164 35649
rect 23848 35640 23900 35692
rect 24400 35640 24452 35692
rect 24952 35683 25004 35692
rect 24952 35649 24961 35683
rect 24961 35649 24995 35683
rect 24995 35649 25004 35683
rect 24952 35640 25004 35649
rect 27160 35708 27212 35760
rect 28080 35708 28132 35760
rect 36360 35776 36412 35828
rect 25688 35683 25740 35692
rect 25688 35649 25697 35683
rect 25697 35649 25731 35683
rect 25731 35649 25740 35683
rect 25688 35640 25740 35649
rect 27712 35640 27764 35692
rect 34520 35640 34572 35692
rect 34704 35683 34756 35692
rect 34704 35649 34713 35683
rect 34713 35649 34747 35683
rect 34747 35649 34756 35683
rect 34704 35640 34756 35649
rect 36544 35640 36596 35692
rect 3240 35572 3292 35624
rect 17224 35479 17276 35488
rect 17224 35445 17233 35479
rect 17233 35445 17267 35479
rect 17267 35445 17276 35479
rect 17224 35436 17276 35445
rect 24584 35572 24636 35624
rect 24860 35615 24912 35624
rect 24860 35581 24869 35615
rect 24869 35581 24903 35615
rect 24903 35581 24912 35615
rect 24860 35572 24912 35581
rect 33784 35572 33836 35624
rect 34612 35572 34664 35624
rect 35440 35572 35492 35624
rect 38108 35615 38160 35624
rect 38108 35581 38117 35615
rect 38117 35581 38151 35615
rect 38151 35581 38160 35615
rect 38108 35572 38160 35581
rect 24308 35504 24360 35556
rect 30656 35504 30708 35556
rect 20168 35436 20220 35488
rect 21272 35479 21324 35488
rect 21272 35445 21281 35479
rect 21281 35445 21315 35479
rect 21315 35445 21324 35479
rect 21272 35436 21324 35445
rect 23756 35436 23808 35488
rect 24768 35436 24820 35488
rect 24860 35436 24912 35488
rect 25872 35436 25924 35488
rect 33232 35479 33284 35488
rect 33232 35445 33241 35479
rect 33241 35445 33275 35479
rect 33275 35445 33284 35479
rect 33232 35436 33284 35445
rect 34796 35436 34848 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 17408 35275 17460 35284
rect 17408 35241 17417 35275
rect 17417 35241 17451 35275
rect 17451 35241 17460 35275
rect 17408 35232 17460 35241
rect 20904 35232 20956 35284
rect 15568 35071 15620 35080
rect 15568 35037 15577 35071
rect 15577 35037 15611 35071
rect 15611 35037 15620 35071
rect 15568 35028 15620 35037
rect 18328 35071 18380 35080
rect 15936 34960 15988 35012
rect 18328 35037 18337 35071
rect 18337 35037 18371 35071
rect 18371 35037 18380 35071
rect 18328 35028 18380 35037
rect 24860 35232 24912 35284
rect 23388 35164 23440 35216
rect 18696 35028 18748 35080
rect 20812 35028 20864 35080
rect 22744 35028 22796 35080
rect 17868 34960 17920 35012
rect 23756 35164 23808 35216
rect 24584 35207 24636 35216
rect 24584 35173 24593 35207
rect 24593 35173 24627 35207
rect 24627 35173 24636 35207
rect 24584 35164 24636 35173
rect 24860 35139 24912 35148
rect 24860 35105 24869 35139
rect 24869 35105 24903 35139
rect 24903 35105 24912 35139
rect 24860 35096 24912 35105
rect 25780 35139 25832 35148
rect 25780 35105 25789 35139
rect 25789 35105 25823 35139
rect 25823 35105 25832 35139
rect 25780 35096 25832 35105
rect 27068 35232 27120 35284
rect 36544 35275 36596 35284
rect 36544 35241 36553 35275
rect 36553 35241 36587 35275
rect 36587 35241 36596 35275
rect 36544 35232 36596 35241
rect 26424 35164 26476 35216
rect 27160 35139 27212 35148
rect 27160 35105 27169 35139
rect 27169 35105 27203 35139
rect 27203 35105 27212 35139
rect 27160 35096 27212 35105
rect 29552 35096 29604 35148
rect 29644 35096 29696 35148
rect 30196 35139 30248 35148
rect 30196 35105 30205 35139
rect 30205 35105 30239 35139
rect 30239 35105 30248 35139
rect 30196 35096 30248 35105
rect 36360 35096 36412 35148
rect 23848 35071 23900 35080
rect 23848 35037 23857 35071
rect 23857 35037 23891 35071
rect 23891 35037 23900 35071
rect 23848 35028 23900 35037
rect 25044 35028 25096 35080
rect 25688 35071 25740 35080
rect 25688 35037 25697 35071
rect 25697 35037 25731 35071
rect 25731 35037 25740 35071
rect 25688 35028 25740 35037
rect 23112 34960 23164 35012
rect 23480 34960 23532 35012
rect 27528 35028 27580 35080
rect 27896 34960 27948 35012
rect 19248 34892 19300 34944
rect 22560 34892 22612 34944
rect 24860 34892 24912 34944
rect 26056 34892 26108 34944
rect 26332 34892 26384 34944
rect 27436 34892 27488 34944
rect 28172 35071 28224 35080
rect 28172 35037 28181 35071
rect 28181 35037 28215 35071
rect 28215 35037 28224 35071
rect 29920 35071 29972 35080
rect 28172 35028 28224 35037
rect 29920 35037 29929 35071
rect 29929 35037 29963 35071
rect 29963 35037 29972 35071
rect 29920 35028 29972 35037
rect 32036 35028 32088 35080
rect 32864 35028 32916 35080
rect 36176 35028 36228 35080
rect 37464 35071 37516 35080
rect 31852 35003 31904 35012
rect 31852 34969 31861 35003
rect 31861 34969 31895 35003
rect 31895 34969 31904 35003
rect 31852 34960 31904 34969
rect 32128 34960 32180 35012
rect 33232 34960 33284 35012
rect 34796 34960 34848 35012
rect 35808 34960 35860 35012
rect 37464 35037 37473 35071
rect 37473 35037 37507 35071
rect 37507 35037 37516 35071
rect 37464 35028 37516 35037
rect 30472 34892 30524 34944
rect 31944 34935 31996 34944
rect 31944 34901 31953 34935
rect 31953 34901 31987 34935
rect 31987 34901 31996 34935
rect 31944 34892 31996 34901
rect 34612 34892 34664 34944
rect 37556 34892 37608 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 15936 34731 15988 34740
rect 15936 34697 15945 34731
rect 15945 34697 15979 34731
rect 15979 34697 15988 34731
rect 15936 34688 15988 34697
rect 18328 34731 18380 34740
rect 18328 34697 18337 34731
rect 18337 34697 18371 34731
rect 18371 34697 18380 34731
rect 18328 34688 18380 34697
rect 20812 34731 20864 34740
rect 20812 34697 20821 34731
rect 20821 34697 20855 34731
rect 20855 34697 20864 34731
rect 20812 34688 20864 34697
rect 22560 34688 22612 34740
rect 23848 34688 23900 34740
rect 17224 34663 17276 34672
rect 17224 34629 17258 34663
rect 17258 34629 17276 34663
rect 17224 34620 17276 34629
rect 16672 34552 16724 34604
rect 19432 34552 19484 34604
rect 21088 34552 21140 34604
rect 21272 34552 21324 34604
rect 21640 34552 21692 34604
rect 22836 34620 22888 34672
rect 26976 34688 27028 34740
rect 22744 34595 22796 34604
rect 22744 34561 22753 34595
rect 22753 34561 22787 34595
rect 22787 34561 22796 34595
rect 23480 34595 23532 34604
rect 22744 34552 22796 34561
rect 15200 34484 15252 34536
rect 15568 34484 15620 34536
rect 16488 34484 16540 34536
rect 20168 34527 20220 34536
rect 20168 34493 20177 34527
rect 20177 34493 20211 34527
rect 20211 34493 20220 34527
rect 20168 34484 20220 34493
rect 22836 34484 22888 34536
rect 23480 34561 23489 34595
rect 23489 34561 23523 34595
rect 23523 34561 23532 34595
rect 23480 34552 23532 34561
rect 23572 34552 23624 34604
rect 24308 34552 24360 34604
rect 24676 34595 24728 34604
rect 24676 34561 24685 34595
rect 24685 34561 24719 34595
rect 24719 34561 24728 34595
rect 24676 34552 24728 34561
rect 24768 34595 24820 34604
rect 24768 34561 24777 34595
rect 24777 34561 24811 34595
rect 24811 34561 24820 34595
rect 25044 34595 25096 34604
rect 24768 34552 24820 34561
rect 25044 34561 25053 34595
rect 25053 34561 25087 34595
rect 25087 34561 25096 34595
rect 26332 34620 26384 34672
rect 25044 34552 25096 34561
rect 24860 34527 24912 34536
rect 24860 34493 24869 34527
rect 24869 34493 24903 34527
rect 24903 34493 24912 34527
rect 24860 34484 24912 34493
rect 24492 34416 24544 34468
rect 26424 34595 26476 34604
rect 26424 34561 26433 34595
rect 26433 34561 26467 34595
rect 26467 34561 26476 34595
rect 26424 34552 26476 34561
rect 26608 34552 26660 34604
rect 27344 34595 27396 34604
rect 27344 34561 27353 34595
rect 27353 34561 27387 34595
rect 27387 34561 27396 34595
rect 27344 34552 27396 34561
rect 27712 34552 27764 34604
rect 28448 34552 28500 34604
rect 29920 34688 29972 34740
rect 33232 34688 33284 34740
rect 34520 34688 34572 34740
rect 37004 34688 37056 34740
rect 32588 34620 32640 34672
rect 34612 34620 34664 34672
rect 35900 34620 35952 34672
rect 30564 34552 30616 34604
rect 34428 34552 34480 34604
rect 35440 34595 35492 34604
rect 35440 34561 35449 34595
rect 35449 34561 35483 34595
rect 35483 34561 35492 34595
rect 35440 34552 35492 34561
rect 27988 34484 28040 34536
rect 28264 34527 28316 34536
rect 28264 34493 28273 34527
rect 28273 34493 28307 34527
rect 28307 34493 28316 34527
rect 28264 34484 28316 34493
rect 29092 34484 29144 34536
rect 26424 34416 26476 34468
rect 28080 34416 28132 34468
rect 29552 34527 29604 34536
rect 29552 34493 29561 34527
rect 29561 34493 29595 34527
rect 29595 34493 29604 34527
rect 29552 34484 29604 34493
rect 32036 34484 32088 34536
rect 33968 34527 34020 34536
rect 33968 34493 33977 34527
rect 33977 34493 34011 34527
rect 34011 34493 34020 34527
rect 33968 34484 34020 34493
rect 36360 34484 36412 34536
rect 36728 34620 36780 34672
rect 37556 34595 37608 34604
rect 37556 34561 37565 34595
rect 37565 34561 37599 34595
rect 37599 34561 37608 34595
rect 37556 34552 37608 34561
rect 18144 34348 18196 34400
rect 25320 34348 25372 34400
rect 26884 34348 26936 34400
rect 34796 34348 34848 34400
rect 36360 34391 36412 34400
rect 36360 34357 36369 34391
rect 36369 34357 36403 34391
rect 36403 34357 36412 34391
rect 36360 34348 36412 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 16672 34187 16724 34196
rect 16672 34153 16681 34187
rect 16681 34153 16715 34187
rect 16715 34153 16724 34187
rect 16672 34144 16724 34153
rect 19432 34187 19484 34196
rect 19432 34153 19441 34187
rect 19441 34153 19475 34187
rect 19475 34153 19484 34187
rect 19432 34144 19484 34153
rect 25688 34144 25740 34196
rect 28172 34144 28224 34196
rect 30564 34187 30616 34196
rect 30564 34153 30573 34187
rect 30573 34153 30607 34187
rect 30607 34153 30616 34187
rect 30564 34144 30616 34153
rect 34704 34187 34756 34196
rect 34704 34153 34713 34187
rect 34713 34153 34747 34187
rect 34747 34153 34756 34187
rect 34704 34144 34756 34153
rect 35900 34144 35952 34196
rect 17868 34119 17920 34128
rect 17868 34085 17877 34119
rect 17877 34085 17911 34119
rect 17911 34085 17920 34119
rect 17868 34076 17920 34085
rect 16856 33983 16908 33992
rect 16856 33949 16865 33983
rect 16865 33949 16899 33983
rect 16899 33949 16908 33983
rect 16856 33940 16908 33949
rect 25044 34008 25096 34060
rect 18144 33983 18196 33992
rect 15108 33915 15160 33924
rect 15108 33881 15142 33915
rect 15142 33881 15160 33915
rect 15108 33872 15160 33881
rect 15200 33872 15252 33924
rect 18144 33949 18153 33983
rect 18153 33949 18187 33983
rect 18187 33949 18196 33983
rect 18144 33940 18196 33949
rect 18328 33940 18380 33992
rect 19248 33983 19300 33992
rect 19248 33949 19257 33983
rect 19257 33949 19291 33983
rect 19291 33949 19300 33983
rect 19248 33940 19300 33949
rect 20168 33940 20220 33992
rect 23020 33940 23072 33992
rect 24492 33983 24544 33992
rect 24492 33949 24501 33983
rect 24501 33949 24535 33983
rect 24535 33949 24544 33983
rect 24492 33940 24544 33949
rect 24952 33940 25004 33992
rect 26792 34008 26844 34060
rect 26884 33983 26936 33992
rect 26884 33949 26893 33983
rect 26893 33949 26927 33983
rect 26927 33949 26936 33983
rect 26884 33940 26936 33949
rect 26976 33983 27028 33992
rect 26976 33949 26985 33983
rect 26985 33949 27019 33983
rect 27019 33949 27028 33983
rect 26976 33940 27028 33949
rect 28080 33983 28132 33992
rect 20904 33872 20956 33924
rect 28080 33949 28089 33983
rect 28089 33949 28123 33983
rect 28123 33949 28132 33983
rect 28080 33940 28132 33949
rect 28264 33983 28316 33992
rect 28264 33949 28273 33983
rect 28273 33949 28307 33983
rect 28307 33949 28316 33983
rect 28264 33940 28316 33949
rect 28448 33940 28500 33992
rect 29092 34008 29144 34060
rect 30656 34076 30708 34128
rect 32956 34076 33008 34128
rect 37740 34144 37792 34196
rect 32128 34051 32180 34060
rect 29552 33940 29604 33992
rect 30472 33940 30524 33992
rect 32128 34017 32137 34051
rect 32137 34017 32171 34051
rect 32171 34017 32180 34051
rect 32128 34008 32180 34017
rect 33784 34051 33836 34060
rect 33784 34017 33793 34051
rect 33793 34017 33827 34051
rect 33827 34017 33836 34051
rect 33784 34008 33836 34017
rect 34520 34008 34572 34060
rect 32220 33940 32272 33992
rect 33692 33983 33744 33992
rect 33692 33949 33701 33983
rect 33701 33949 33735 33983
rect 33735 33949 33744 33983
rect 33692 33940 33744 33949
rect 35808 34008 35860 34060
rect 36176 34008 36228 34060
rect 18052 33847 18104 33856
rect 18052 33813 18061 33847
rect 18061 33813 18095 33847
rect 18095 33813 18104 33847
rect 18052 33804 18104 33813
rect 18420 33847 18472 33856
rect 18420 33813 18429 33847
rect 18429 33813 18463 33847
rect 18463 33813 18472 33847
rect 18420 33804 18472 33813
rect 20076 33804 20128 33856
rect 28540 33804 28592 33856
rect 29828 33804 29880 33856
rect 31944 33804 31996 33856
rect 33324 33804 33376 33856
rect 33508 33847 33560 33856
rect 33508 33813 33517 33847
rect 33517 33813 33551 33847
rect 33551 33813 33560 33847
rect 33508 33804 33560 33813
rect 34612 33872 34664 33924
rect 37464 33940 37516 33992
rect 36268 33915 36320 33924
rect 36268 33881 36277 33915
rect 36277 33881 36311 33915
rect 36311 33881 36320 33915
rect 36268 33872 36320 33881
rect 37004 33915 37056 33924
rect 37004 33881 37038 33915
rect 37038 33881 37056 33915
rect 37004 33872 37056 33881
rect 37556 33804 37608 33856
rect 38108 33847 38160 33856
rect 38108 33813 38117 33847
rect 38117 33813 38151 33847
rect 38151 33813 38160 33847
rect 38108 33804 38160 33813
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 15108 33600 15160 33652
rect 17960 33600 18012 33652
rect 27344 33600 27396 33652
rect 30656 33600 30708 33652
rect 33692 33600 33744 33652
rect 18328 33532 18380 33584
rect 21088 33532 21140 33584
rect 27528 33575 27580 33584
rect 15384 33507 15436 33516
rect 15384 33473 15393 33507
rect 15393 33473 15427 33507
rect 15427 33473 15436 33507
rect 15384 33464 15436 33473
rect 17868 33464 17920 33516
rect 20996 33507 21048 33516
rect 20996 33473 21005 33507
rect 21005 33473 21039 33507
rect 21039 33473 21048 33507
rect 20996 33464 21048 33473
rect 23020 33464 23072 33516
rect 25320 33507 25372 33516
rect 25320 33473 25354 33507
rect 25354 33473 25372 33507
rect 25320 33464 25372 33473
rect 18144 33439 18196 33448
rect 18144 33405 18153 33439
rect 18153 33405 18187 33439
rect 18187 33405 18196 33439
rect 18144 33396 18196 33405
rect 27528 33541 27537 33575
rect 27537 33541 27571 33575
rect 27571 33541 27580 33575
rect 27528 33532 27580 33541
rect 29644 33575 29696 33584
rect 29644 33541 29653 33575
rect 29653 33541 29687 33575
rect 29687 33541 29696 33575
rect 29644 33532 29696 33541
rect 36268 33532 36320 33584
rect 27436 33464 27488 33516
rect 30380 33507 30432 33516
rect 30380 33473 30389 33507
rect 30389 33473 30423 33507
rect 30423 33473 30432 33507
rect 30380 33464 30432 33473
rect 34428 33507 34480 33516
rect 34428 33473 34437 33507
rect 34437 33473 34471 33507
rect 34471 33473 34480 33507
rect 34428 33464 34480 33473
rect 34796 33464 34848 33516
rect 37280 33464 37332 33516
rect 38108 33532 38160 33584
rect 37556 33507 37608 33516
rect 37556 33473 37565 33507
rect 37565 33473 37599 33507
rect 37599 33473 37608 33507
rect 37556 33464 37608 33473
rect 37740 33507 37792 33516
rect 37740 33473 37749 33507
rect 37749 33473 37783 33507
rect 37783 33473 37792 33507
rect 37740 33464 37792 33473
rect 31300 33396 31352 33448
rect 21824 33328 21876 33380
rect 23112 33328 23164 33380
rect 18052 33303 18104 33312
rect 18052 33269 18061 33303
rect 18061 33269 18095 33303
rect 18095 33269 18104 33303
rect 18052 33260 18104 33269
rect 22008 33303 22060 33312
rect 22008 33269 22017 33303
rect 22017 33269 22051 33303
rect 22051 33269 22060 33303
rect 22008 33260 22060 33269
rect 22836 33260 22888 33312
rect 33968 33328 34020 33380
rect 34520 33328 34572 33380
rect 26424 33303 26476 33312
rect 26424 33269 26433 33303
rect 26433 33269 26467 33303
rect 26467 33269 26476 33303
rect 26424 33260 26476 33269
rect 26976 33260 27028 33312
rect 29828 33260 29880 33312
rect 36452 33303 36504 33312
rect 36452 33269 36461 33303
rect 36461 33269 36495 33303
rect 36495 33269 36504 33303
rect 36452 33260 36504 33269
rect 37464 33303 37516 33312
rect 37464 33269 37473 33303
rect 37473 33269 37507 33303
rect 37507 33269 37516 33303
rect 37464 33260 37516 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 15384 33099 15436 33108
rect 15384 33065 15393 33099
rect 15393 33065 15427 33099
rect 15427 33065 15436 33099
rect 15384 33056 15436 33065
rect 16856 33056 16908 33108
rect 32404 33056 32456 33108
rect 33140 33056 33192 33108
rect 37556 33099 37608 33108
rect 37556 33065 37565 33099
rect 37565 33065 37599 33099
rect 37599 33065 37608 33099
rect 37556 33056 37608 33065
rect 15568 32895 15620 32904
rect 15568 32861 15577 32895
rect 15577 32861 15611 32895
rect 15611 32861 15620 32895
rect 15568 32852 15620 32861
rect 15660 32895 15712 32904
rect 15660 32861 15669 32895
rect 15669 32861 15703 32895
rect 15703 32861 15712 32895
rect 18604 32920 18656 32972
rect 20996 32920 21048 32972
rect 34520 32920 34572 32972
rect 35808 32920 35860 32972
rect 36176 32963 36228 32972
rect 36176 32929 36185 32963
rect 36185 32929 36219 32963
rect 36219 32929 36228 32963
rect 36176 32920 36228 32929
rect 15660 32852 15712 32861
rect 17960 32895 18012 32904
rect 17960 32861 17969 32895
rect 17969 32861 18003 32895
rect 18003 32861 18012 32895
rect 17960 32852 18012 32861
rect 23664 32852 23716 32904
rect 30380 32852 30432 32904
rect 32220 32895 32272 32904
rect 16948 32784 17000 32836
rect 32220 32861 32229 32895
rect 32229 32861 32263 32895
rect 32263 32861 32272 32895
rect 32220 32852 32272 32861
rect 36452 32895 36504 32904
rect 36452 32861 36486 32895
rect 36486 32861 36504 32895
rect 36452 32852 36504 32861
rect 33232 32784 33284 32836
rect 18512 32716 18564 32768
rect 23664 32759 23716 32768
rect 23664 32725 23673 32759
rect 23673 32725 23707 32759
rect 23707 32725 23716 32759
rect 23664 32716 23716 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 15660 32555 15712 32564
rect 15660 32521 15669 32555
rect 15669 32521 15703 32555
rect 15703 32521 15712 32555
rect 15660 32512 15712 32521
rect 16672 32512 16724 32564
rect 23572 32512 23624 32564
rect 30932 32512 30984 32564
rect 37280 32555 37332 32564
rect 37280 32521 37289 32555
rect 37289 32521 37323 32555
rect 37323 32521 37332 32555
rect 37280 32512 37332 32521
rect 15200 32444 15252 32496
rect 14556 32419 14608 32428
rect 14556 32385 14590 32419
rect 14590 32385 14608 32419
rect 14556 32376 14608 32385
rect 16764 32376 16816 32428
rect 17040 32419 17092 32428
rect 17040 32385 17049 32419
rect 17049 32385 17083 32419
rect 17083 32385 17092 32419
rect 17040 32376 17092 32385
rect 18328 32376 18380 32428
rect 20996 32376 21048 32428
rect 23020 32444 23072 32496
rect 27528 32444 27580 32496
rect 30380 32444 30432 32496
rect 30472 32487 30524 32496
rect 30472 32453 30497 32487
rect 30497 32453 30524 32487
rect 31300 32487 31352 32496
rect 30472 32444 30524 32453
rect 31300 32453 31309 32487
rect 31309 32453 31343 32487
rect 31343 32453 31352 32487
rect 31300 32444 31352 32453
rect 32220 32444 32272 32496
rect 33508 32444 33560 32496
rect 35808 32444 35860 32496
rect 23204 32376 23256 32428
rect 20628 32351 20680 32360
rect 16580 32240 16632 32292
rect 20628 32317 20637 32351
rect 20637 32317 20671 32351
rect 20671 32317 20680 32351
rect 20628 32308 20680 32317
rect 24860 32376 24912 32428
rect 25412 32419 25464 32428
rect 25412 32385 25421 32419
rect 25421 32385 25455 32419
rect 25455 32385 25464 32419
rect 25412 32376 25464 32385
rect 25872 32376 25924 32428
rect 25780 32308 25832 32360
rect 27896 32240 27948 32292
rect 28908 32376 28960 32428
rect 32496 32419 32548 32428
rect 32496 32385 32505 32419
rect 32505 32385 32539 32419
rect 32539 32385 32548 32419
rect 32496 32376 32548 32385
rect 36268 32419 36320 32428
rect 36268 32385 36277 32419
rect 36277 32385 36311 32419
rect 36311 32385 36320 32419
rect 36268 32376 36320 32385
rect 37740 32376 37792 32428
rect 28448 32308 28500 32360
rect 29828 32308 29880 32360
rect 32036 32308 32088 32360
rect 28264 32240 28316 32292
rect 28632 32240 28684 32292
rect 18236 32172 18288 32224
rect 20260 32215 20312 32224
rect 20260 32181 20269 32215
rect 20269 32181 20303 32215
rect 20303 32181 20312 32215
rect 20260 32172 20312 32181
rect 23940 32215 23992 32224
rect 23940 32181 23949 32215
rect 23949 32181 23983 32215
rect 23983 32181 23992 32215
rect 23940 32172 23992 32181
rect 27160 32172 27212 32224
rect 28356 32172 28408 32224
rect 30380 32172 30432 32224
rect 33232 32172 33284 32224
rect 35440 32215 35492 32224
rect 35440 32181 35449 32215
rect 35449 32181 35483 32215
rect 35483 32181 35492 32215
rect 35440 32172 35492 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 14556 31968 14608 32020
rect 16764 32011 16816 32020
rect 16764 31977 16773 32011
rect 16773 31977 16807 32011
rect 16807 31977 16816 32011
rect 16764 31968 16816 31977
rect 16948 32011 17000 32020
rect 16948 31977 16957 32011
rect 16957 31977 16991 32011
rect 16991 31977 17000 32011
rect 16948 31968 17000 31977
rect 18328 31968 18380 32020
rect 18604 31968 18656 32020
rect 22008 31968 22060 32020
rect 23204 32011 23256 32020
rect 23204 31977 23213 32011
rect 23213 31977 23247 32011
rect 23247 31977 23256 32011
rect 23204 31968 23256 31977
rect 26240 31968 26292 32020
rect 30748 31968 30800 32020
rect 30932 32011 30984 32020
rect 30932 31977 30941 32011
rect 30941 31977 30975 32011
rect 30975 31977 30984 32011
rect 30932 31968 30984 31977
rect 15568 31807 15620 31816
rect 15568 31773 15577 31807
rect 15577 31773 15611 31807
rect 15611 31773 15620 31807
rect 15568 31764 15620 31773
rect 17040 31900 17092 31952
rect 16672 31875 16724 31884
rect 16672 31841 16681 31875
rect 16681 31841 16715 31875
rect 16715 31841 16724 31875
rect 16672 31832 16724 31841
rect 18236 31807 18288 31816
rect 16672 31696 16724 31748
rect 18236 31773 18245 31807
rect 18245 31773 18279 31807
rect 18279 31773 18288 31807
rect 18236 31764 18288 31773
rect 18420 31832 18472 31884
rect 18696 31875 18748 31884
rect 18696 31841 18705 31875
rect 18705 31841 18739 31875
rect 18739 31841 18748 31875
rect 18696 31832 18748 31841
rect 18512 31807 18564 31816
rect 18512 31773 18547 31807
rect 18547 31773 18564 31807
rect 20720 31900 20772 31952
rect 21272 31900 21324 31952
rect 22744 31900 22796 31952
rect 23020 31900 23072 31952
rect 27344 31900 27396 31952
rect 32496 31900 32548 31952
rect 34428 31968 34480 32020
rect 20628 31875 20680 31884
rect 20628 31841 20637 31875
rect 20637 31841 20671 31875
rect 20671 31841 20680 31875
rect 20628 31832 20680 31841
rect 20996 31832 21048 31884
rect 18512 31764 18564 31773
rect 20260 31764 20312 31816
rect 23388 31832 23440 31884
rect 30380 31832 30432 31884
rect 23940 31764 23992 31816
rect 24584 31807 24636 31816
rect 23664 31696 23716 31748
rect 24584 31773 24593 31807
rect 24593 31773 24627 31807
rect 24627 31773 24636 31807
rect 24584 31764 24636 31773
rect 25044 31764 25096 31816
rect 27344 31807 27396 31816
rect 27344 31773 27353 31807
rect 27353 31773 27387 31807
rect 27387 31773 27396 31807
rect 27344 31764 27396 31773
rect 28908 31764 28960 31816
rect 29552 31807 29604 31816
rect 29552 31773 29561 31807
rect 29561 31773 29595 31807
rect 29595 31773 29604 31807
rect 29552 31764 29604 31773
rect 29828 31773 29837 31794
rect 29837 31773 29871 31794
rect 29871 31773 29880 31794
rect 29828 31742 29880 31773
rect 29920 31807 29972 31816
rect 29920 31773 29929 31807
rect 29929 31773 29963 31807
rect 29963 31773 29972 31807
rect 29920 31764 29972 31773
rect 30196 31764 30248 31816
rect 31300 31764 31352 31816
rect 31760 31764 31812 31816
rect 35348 31900 35400 31952
rect 37464 31832 37516 31884
rect 38108 31875 38160 31884
rect 38108 31841 38117 31875
rect 38117 31841 38151 31875
rect 38151 31841 38160 31875
rect 38108 31832 38160 31841
rect 33232 31764 33284 31816
rect 26056 31628 26108 31680
rect 29460 31628 29512 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 10968 31424 11020 31476
rect 18696 31399 18748 31408
rect 15568 31331 15620 31340
rect 15568 31297 15574 31331
rect 15574 31297 15608 31331
rect 15608 31297 15620 31331
rect 15568 31288 15620 31297
rect 16764 31288 16816 31340
rect 18696 31365 18730 31399
rect 18730 31365 18748 31399
rect 18696 31356 18748 31365
rect 20076 31356 20128 31408
rect 20628 31288 20680 31340
rect 21272 31356 21324 31408
rect 23020 31399 23072 31408
rect 23020 31365 23054 31399
rect 23054 31365 23072 31399
rect 23020 31356 23072 31365
rect 21824 31288 21876 31340
rect 16672 31263 16724 31272
rect 16672 31229 16681 31263
rect 16681 31229 16715 31263
rect 16715 31229 16724 31263
rect 16672 31220 16724 31229
rect 18420 31263 18472 31272
rect 18420 31229 18429 31263
rect 18429 31229 18463 31263
rect 18463 31229 18472 31263
rect 18420 31220 18472 31229
rect 20812 31263 20864 31272
rect 20812 31229 20821 31263
rect 20821 31229 20855 31263
rect 20855 31229 20864 31263
rect 20812 31220 20864 31229
rect 22468 31220 22520 31272
rect 24768 31288 24820 31340
rect 25228 31424 25280 31476
rect 25412 31467 25464 31476
rect 25412 31433 25421 31467
rect 25421 31433 25455 31467
rect 25455 31433 25464 31467
rect 25412 31424 25464 31433
rect 25780 31424 25832 31476
rect 26056 31424 26108 31476
rect 26056 31331 26108 31340
rect 26056 31297 26065 31331
rect 26065 31297 26099 31331
rect 26099 31297 26108 31331
rect 26056 31288 26108 31297
rect 26332 31288 26384 31340
rect 29276 31424 29328 31476
rect 28540 31399 28592 31408
rect 28540 31365 28558 31399
rect 28558 31365 28592 31399
rect 28540 31356 28592 31365
rect 27160 31288 27212 31340
rect 28080 31288 28132 31340
rect 29460 31331 29512 31340
rect 29460 31297 29469 31331
rect 29469 31297 29503 31331
rect 29503 31297 29512 31331
rect 29460 31288 29512 31297
rect 30012 31424 30064 31476
rect 30380 31424 30432 31476
rect 30932 31424 30984 31476
rect 37464 31424 37516 31476
rect 29736 31331 29788 31340
rect 29736 31297 29745 31331
rect 29745 31297 29779 31331
rect 29779 31297 29788 31331
rect 29736 31288 29788 31297
rect 31300 31288 31352 31340
rect 31668 31288 31720 31340
rect 32404 31331 32456 31340
rect 32404 31297 32438 31331
rect 32438 31297 32456 31331
rect 32404 31288 32456 31297
rect 35440 31356 35492 31408
rect 37556 31288 37608 31340
rect 14280 31084 14332 31136
rect 17684 31127 17736 31136
rect 17684 31093 17693 31127
rect 17693 31093 17727 31127
rect 17727 31093 17736 31127
rect 17684 31084 17736 31093
rect 21180 31127 21232 31136
rect 21180 31093 21189 31127
rect 21189 31093 21223 31127
rect 21223 31093 21232 31127
rect 21180 31084 21232 31093
rect 25504 31084 25556 31136
rect 27436 31127 27488 31136
rect 27436 31093 27445 31127
rect 27445 31093 27479 31127
rect 27479 31093 27488 31127
rect 27436 31084 27488 31093
rect 32036 31220 32088 31272
rect 34060 31220 34112 31272
rect 33784 31084 33836 31136
rect 37740 31152 37792 31204
rect 37556 31084 37608 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 2136 30880 2188 30932
rect 25872 30923 25924 30932
rect 16672 30812 16724 30864
rect 17040 30812 17092 30864
rect 20628 30812 20680 30864
rect 21272 30744 21324 30796
rect 25872 30889 25881 30923
rect 25881 30889 25915 30923
rect 25915 30889 25924 30923
rect 25872 30880 25924 30889
rect 27528 30923 27580 30932
rect 27528 30889 27537 30923
rect 27537 30889 27571 30923
rect 27571 30889 27580 30923
rect 27528 30880 27580 30889
rect 24492 30812 24544 30864
rect 29460 30880 29512 30932
rect 29736 30880 29788 30932
rect 28632 30812 28684 30864
rect 32404 30787 32456 30796
rect 32404 30753 32413 30787
rect 32413 30753 32447 30787
rect 32447 30753 32456 30787
rect 32404 30744 32456 30753
rect 37188 30787 37240 30796
rect 37188 30753 37197 30787
rect 37197 30753 37231 30787
rect 37231 30753 37240 30787
rect 37188 30744 37240 30753
rect 37280 30744 37332 30796
rect 37924 30744 37976 30796
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 18052 30676 18104 30728
rect 18420 30676 18472 30728
rect 20076 30719 20128 30728
rect 20076 30685 20085 30719
rect 20085 30685 20119 30719
rect 20119 30685 20128 30719
rect 20076 30676 20128 30685
rect 20812 30676 20864 30728
rect 21824 30719 21876 30728
rect 21824 30685 21833 30719
rect 21833 30685 21867 30719
rect 21867 30685 21876 30719
rect 21824 30676 21876 30685
rect 22836 30676 22888 30728
rect 24768 30719 24820 30728
rect 24768 30685 24777 30719
rect 24777 30685 24811 30719
rect 24811 30685 24820 30719
rect 24768 30676 24820 30685
rect 25504 30719 25556 30728
rect 17684 30608 17736 30660
rect 20904 30608 20956 30660
rect 24492 30608 24544 30660
rect 25504 30685 25513 30719
rect 25513 30685 25547 30719
rect 25547 30685 25556 30719
rect 25504 30676 25556 30685
rect 26976 30676 27028 30728
rect 26424 30608 26476 30660
rect 27436 30676 27488 30728
rect 28080 30719 28132 30728
rect 28080 30685 28089 30719
rect 28089 30685 28123 30719
rect 28123 30685 28132 30719
rect 28080 30676 28132 30685
rect 28356 30719 28408 30728
rect 28356 30685 28365 30719
rect 28365 30685 28399 30719
rect 28399 30685 28408 30719
rect 28356 30676 28408 30685
rect 30932 30676 30984 30728
rect 31852 30719 31904 30728
rect 31852 30685 31861 30719
rect 31861 30685 31895 30719
rect 31895 30685 31904 30719
rect 31852 30676 31904 30685
rect 38200 30676 38252 30728
rect 37924 30651 37976 30660
rect 37924 30617 37933 30651
rect 37933 30617 37967 30651
rect 37967 30617 37976 30651
rect 37924 30608 37976 30617
rect 21088 30540 21140 30592
rect 21916 30540 21968 30592
rect 23296 30540 23348 30592
rect 26608 30540 26660 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 21088 30336 21140 30388
rect 22008 30336 22060 30388
rect 27528 30379 27580 30388
rect 27528 30345 27537 30379
rect 27537 30345 27571 30379
rect 27571 30345 27580 30379
rect 27528 30336 27580 30345
rect 14924 30243 14976 30252
rect 14924 30209 14933 30243
rect 14933 30209 14967 30243
rect 14967 30209 14976 30243
rect 14924 30200 14976 30209
rect 18604 30243 18656 30252
rect 18604 30209 18613 30243
rect 18613 30209 18647 30243
rect 18647 30209 18656 30243
rect 18604 30200 18656 30209
rect 20904 30243 20956 30252
rect 15384 30175 15436 30184
rect 15384 30141 15393 30175
rect 15393 30141 15427 30175
rect 15427 30141 15436 30175
rect 15384 30132 15436 30141
rect 18604 29996 18656 30048
rect 20904 30209 20913 30243
rect 20913 30209 20947 30243
rect 20947 30209 20956 30243
rect 20904 30200 20956 30209
rect 21088 30243 21140 30252
rect 21088 30209 21097 30243
rect 21097 30209 21131 30243
rect 21131 30209 21140 30243
rect 21088 30200 21140 30209
rect 21548 30200 21600 30252
rect 21916 30200 21968 30252
rect 22100 30243 22152 30252
rect 22100 30209 22109 30243
rect 22109 30209 22143 30243
rect 22143 30209 22152 30243
rect 22100 30200 22152 30209
rect 20996 30132 21048 30184
rect 21180 30132 21232 30184
rect 22192 30132 22244 30184
rect 22376 30243 22428 30252
rect 22376 30209 22385 30243
rect 22385 30209 22419 30243
rect 22419 30209 22428 30243
rect 22376 30200 22428 30209
rect 26332 30268 26384 30320
rect 28908 30311 28960 30320
rect 24584 30200 24636 30252
rect 25044 30243 25096 30252
rect 25044 30209 25053 30243
rect 25053 30209 25087 30243
rect 25087 30209 25096 30243
rect 25044 30200 25096 30209
rect 28264 30200 28316 30252
rect 28908 30277 28917 30311
rect 28917 30277 28951 30311
rect 28951 30277 28960 30311
rect 28908 30268 28960 30277
rect 30564 30268 30616 30320
rect 31300 30336 31352 30388
rect 37924 30336 37976 30388
rect 31484 30268 31536 30320
rect 33324 30268 33376 30320
rect 34428 30268 34480 30320
rect 28816 30243 28868 30252
rect 28816 30209 28825 30243
rect 28825 30209 28859 30243
rect 28859 30209 28868 30243
rect 28816 30200 28868 30209
rect 29000 30200 29052 30252
rect 29644 30243 29696 30252
rect 29644 30209 29653 30243
rect 29653 30209 29687 30243
rect 29687 30209 29696 30243
rect 29644 30200 29696 30209
rect 34060 30243 34112 30252
rect 34060 30209 34069 30243
rect 34069 30209 34103 30243
rect 34103 30209 34112 30243
rect 34060 30200 34112 30209
rect 37280 30200 37332 30252
rect 37464 30200 37516 30252
rect 20904 30064 20956 30116
rect 21364 30064 21416 30116
rect 27896 30064 27948 30116
rect 21272 30039 21324 30048
rect 21272 30005 21281 30039
rect 21281 30005 21315 30039
rect 21315 30005 21324 30039
rect 21272 29996 21324 30005
rect 21824 30039 21876 30048
rect 21824 30005 21833 30039
rect 21833 30005 21867 30039
rect 21867 30005 21876 30039
rect 21824 29996 21876 30005
rect 29460 30039 29512 30048
rect 29460 30005 29469 30039
rect 29469 30005 29503 30039
rect 29503 30005 29512 30039
rect 29460 29996 29512 30005
rect 31576 30064 31628 30116
rect 31760 30064 31812 30116
rect 33232 30064 33284 30116
rect 30380 29996 30432 30048
rect 31668 29996 31720 30048
rect 33692 29996 33744 30048
rect 35440 30039 35492 30048
rect 35440 30005 35449 30039
rect 35449 30005 35483 30039
rect 35483 30005 35492 30039
rect 35440 29996 35492 30005
rect 36268 29996 36320 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 20996 29792 21048 29844
rect 15660 29699 15712 29708
rect 15660 29665 15669 29699
rect 15669 29665 15703 29699
rect 15703 29665 15712 29699
rect 15660 29656 15712 29665
rect 18604 29656 18656 29708
rect 21364 29724 21416 29776
rect 22376 29724 22428 29776
rect 22836 29724 22888 29776
rect 21640 29699 21692 29708
rect 21640 29665 21649 29699
rect 21649 29665 21683 29699
rect 21683 29665 21692 29699
rect 21640 29656 21692 29665
rect 1676 29588 1728 29640
rect 14188 29631 14240 29640
rect 14188 29597 14197 29631
rect 14197 29597 14231 29631
rect 14231 29597 14240 29631
rect 14188 29588 14240 29597
rect 14924 29588 14976 29640
rect 20812 29631 20864 29640
rect 20812 29597 20821 29631
rect 20821 29597 20855 29631
rect 20855 29597 20864 29631
rect 20812 29588 20864 29597
rect 20904 29631 20956 29640
rect 20904 29597 20913 29631
rect 20913 29597 20947 29631
rect 20947 29597 20956 29631
rect 20904 29588 20956 29597
rect 21088 29588 21140 29640
rect 22192 29656 22244 29708
rect 25504 29792 25556 29844
rect 26056 29835 26108 29844
rect 26056 29801 26065 29835
rect 26065 29801 26099 29835
rect 26099 29801 26108 29835
rect 26056 29792 26108 29801
rect 26976 29835 27028 29844
rect 26976 29801 26985 29835
rect 26985 29801 27019 29835
rect 27019 29801 27028 29835
rect 26976 29792 27028 29801
rect 29000 29792 29052 29844
rect 30932 29835 30984 29844
rect 27160 29656 27212 29708
rect 22008 29631 22060 29640
rect 22008 29597 22017 29631
rect 22017 29597 22051 29631
rect 22051 29597 22060 29631
rect 22008 29588 22060 29597
rect 23112 29631 23164 29640
rect 15660 29520 15712 29572
rect 14372 29495 14424 29504
rect 14372 29461 14381 29495
rect 14381 29461 14415 29495
rect 14415 29461 14424 29495
rect 14372 29452 14424 29461
rect 20628 29495 20680 29504
rect 20628 29461 20637 29495
rect 20637 29461 20671 29495
rect 20671 29461 20680 29495
rect 20628 29452 20680 29461
rect 21548 29520 21600 29572
rect 23112 29597 23121 29631
rect 23121 29597 23155 29631
rect 23155 29597 23164 29631
rect 23112 29588 23164 29597
rect 25504 29631 25556 29640
rect 25504 29597 25513 29631
rect 25513 29597 25547 29631
rect 25547 29597 25556 29631
rect 25504 29588 25556 29597
rect 25964 29631 26016 29640
rect 25964 29597 25973 29631
rect 25973 29597 26007 29631
rect 26007 29597 26016 29631
rect 25964 29588 26016 29597
rect 26884 29631 26936 29640
rect 26884 29597 26893 29631
rect 26893 29597 26927 29631
rect 26927 29597 26936 29631
rect 26884 29588 26936 29597
rect 28908 29631 28960 29640
rect 28908 29597 28917 29631
rect 28917 29597 28951 29631
rect 28951 29597 28960 29631
rect 28908 29588 28960 29597
rect 29276 29588 29328 29640
rect 30932 29801 30941 29835
rect 30941 29801 30975 29835
rect 30975 29801 30984 29835
rect 30932 29792 30984 29801
rect 30656 29724 30708 29776
rect 33324 29724 33376 29776
rect 34796 29724 34848 29776
rect 33784 29699 33836 29708
rect 33784 29665 33793 29699
rect 33793 29665 33827 29699
rect 33827 29665 33836 29699
rect 33784 29656 33836 29665
rect 30380 29588 30432 29640
rect 31668 29631 31720 29640
rect 31668 29597 31677 29631
rect 31677 29597 31711 29631
rect 31711 29597 31720 29631
rect 31668 29588 31720 29597
rect 34612 29588 34664 29640
rect 35440 29656 35492 29708
rect 36268 29699 36320 29708
rect 36268 29665 36277 29699
rect 36277 29665 36311 29699
rect 36311 29665 36320 29699
rect 36268 29656 36320 29665
rect 38108 29699 38160 29708
rect 38108 29665 38117 29699
rect 38117 29665 38151 29699
rect 38151 29665 38160 29699
rect 38108 29656 38160 29665
rect 29368 29520 29420 29572
rect 29460 29520 29512 29572
rect 30840 29520 30892 29572
rect 33232 29520 33284 29572
rect 34428 29520 34480 29572
rect 37372 29520 37424 29572
rect 23296 29495 23348 29504
rect 23296 29461 23305 29495
rect 23305 29461 23339 29495
rect 23339 29461 23348 29495
rect 23296 29452 23348 29461
rect 24860 29452 24912 29504
rect 31208 29452 31260 29504
rect 31300 29452 31352 29504
rect 33416 29452 33468 29504
rect 34520 29452 34572 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 24860 29248 24912 29300
rect 25412 29248 25464 29300
rect 25964 29248 26016 29300
rect 26884 29248 26936 29300
rect 29644 29291 29696 29300
rect 29644 29257 29653 29291
rect 29653 29257 29687 29291
rect 29687 29257 29696 29291
rect 29644 29248 29696 29257
rect 30564 29248 30616 29300
rect 1676 29155 1728 29164
rect 1676 29121 1685 29155
rect 1685 29121 1719 29155
rect 1719 29121 1728 29155
rect 1676 29112 1728 29121
rect 14096 29155 14148 29164
rect 14096 29121 14105 29155
rect 14105 29121 14139 29155
rect 14139 29121 14148 29155
rect 14372 29155 14424 29164
rect 14096 29112 14148 29121
rect 14372 29121 14381 29155
rect 14381 29121 14415 29155
rect 14415 29121 14424 29155
rect 14924 29155 14976 29164
rect 14372 29112 14424 29121
rect 14924 29121 14933 29155
rect 14933 29121 14967 29155
rect 14967 29121 14976 29155
rect 14924 29112 14976 29121
rect 18052 29112 18104 29164
rect 18236 29155 18288 29164
rect 18236 29121 18270 29155
rect 18270 29121 18288 29155
rect 22468 29155 22520 29164
rect 18236 29112 18288 29121
rect 1860 29087 1912 29096
rect 1860 29053 1869 29087
rect 1869 29053 1903 29087
rect 1903 29053 1912 29087
rect 1860 29044 1912 29053
rect 2780 29087 2832 29096
rect 2780 29053 2789 29087
rect 2789 29053 2823 29087
rect 2823 29053 2832 29087
rect 2780 29044 2832 29053
rect 15660 29087 15712 29096
rect 15660 29053 15669 29087
rect 15669 29053 15703 29087
rect 15703 29053 15712 29087
rect 15660 29044 15712 29053
rect 18144 28908 18196 28960
rect 19340 28985 19349 29006
rect 19349 28985 19383 29006
rect 19383 28985 19392 29006
rect 19340 28954 19392 28985
rect 19432 28908 19484 28960
rect 22468 29121 22477 29155
rect 22477 29121 22511 29155
rect 22511 29121 22520 29155
rect 22468 29112 22520 29121
rect 22744 29155 22796 29164
rect 22744 29121 22778 29155
rect 22778 29121 22796 29155
rect 22744 29112 22796 29121
rect 25504 29180 25556 29232
rect 25320 29112 25372 29164
rect 28724 29180 28776 29232
rect 28908 29180 28960 29232
rect 31668 29248 31720 29300
rect 37372 29291 37424 29300
rect 37372 29257 37381 29291
rect 37381 29257 37415 29291
rect 37415 29257 37424 29291
rect 37372 29248 37424 29257
rect 27620 29112 27672 29164
rect 30656 29155 30708 29164
rect 22836 28908 22888 28960
rect 30656 29121 30665 29155
rect 30665 29121 30699 29155
rect 30699 29121 30708 29155
rect 30656 29112 30708 29121
rect 35808 29180 35860 29232
rect 31300 29112 31352 29164
rect 29276 29087 29328 29096
rect 29276 29053 29285 29087
rect 29285 29053 29319 29087
rect 29319 29053 29328 29087
rect 29276 29044 29328 29053
rect 31208 29044 31260 29096
rect 33784 29112 33836 29164
rect 34428 29155 34480 29164
rect 34428 29121 34437 29155
rect 34437 29121 34471 29155
rect 34471 29121 34480 29155
rect 34428 29112 34480 29121
rect 34612 29155 34664 29164
rect 34612 29121 34621 29155
rect 34621 29121 34655 29155
rect 34655 29121 34664 29155
rect 34612 29112 34664 29121
rect 35624 29112 35676 29164
rect 37280 29155 37332 29164
rect 37280 29121 37289 29155
rect 37289 29121 37323 29155
rect 37323 29121 37332 29155
rect 37280 29112 37332 29121
rect 38200 29112 38252 29164
rect 31944 29044 31996 29096
rect 30380 28976 30432 29028
rect 30656 28976 30708 29028
rect 25136 28951 25188 28960
rect 25136 28917 25145 28951
rect 25145 28917 25179 28951
rect 25179 28917 25188 28951
rect 25136 28908 25188 28917
rect 30932 28908 30984 28960
rect 31852 28908 31904 28960
rect 34612 28951 34664 28960
rect 34612 28917 34621 28951
rect 34621 28917 34655 28951
rect 34655 28917 34664 28951
rect 34612 28908 34664 28917
rect 35808 28951 35860 28960
rect 35808 28917 35817 28951
rect 35817 28917 35851 28951
rect 35851 28917 35860 28951
rect 35808 28908 35860 28917
rect 36728 28951 36780 28960
rect 36728 28917 36737 28951
rect 36737 28917 36771 28951
rect 36771 28917 36780 28951
rect 36728 28908 36780 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 1860 28704 1912 28756
rect 15936 28704 15988 28756
rect 18236 28704 18288 28756
rect 22744 28704 22796 28756
rect 20444 28636 20496 28688
rect 25504 28704 25556 28756
rect 27620 28747 27672 28756
rect 27620 28713 27629 28747
rect 27629 28713 27663 28747
rect 27663 28713 27672 28747
rect 27620 28704 27672 28713
rect 28264 28704 28316 28756
rect 28908 28704 28960 28756
rect 30932 28636 30984 28688
rect 31300 28636 31352 28688
rect 31576 28636 31628 28688
rect 18052 28568 18104 28620
rect 19432 28568 19484 28620
rect 22468 28568 22520 28620
rect 23480 28568 23532 28620
rect 2320 28543 2372 28552
rect 2320 28509 2329 28543
rect 2329 28509 2363 28543
rect 2363 28509 2372 28543
rect 2320 28500 2372 28509
rect 15292 28543 15344 28552
rect 15292 28509 15301 28543
rect 15301 28509 15335 28543
rect 15335 28509 15344 28543
rect 15292 28500 15344 28509
rect 18144 28500 18196 28552
rect 4804 28432 4856 28484
rect 9588 28432 9640 28484
rect 14648 28475 14700 28484
rect 14648 28441 14657 28475
rect 14657 28441 14691 28475
rect 14691 28441 14700 28475
rect 14648 28432 14700 28441
rect 17316 28432 17368 28484
rect 18512 28543 18564 28552
rect 18512 28509 18526 28543
rect 18526 28509 18560 28543
rect 18560 28509 18564 28543
rect 18512 28500 18564 28509
rect 18696 28543 18748 28552
rect 18696 28509 18705 28543
rect 18705 28509 18739 28543
rect 18739 28509 18748 28543
rect 18696 28500 18748 28509
rect 21456 28500 21508 28552
rect 22836 28500 22888 28552
rect 23020 28543 23072 28552
rect 23020 28509 23029 28543
rect 23029 28509 23063 28543
rect 23063 28509 23072 28543
rect 23020 28500 23072 28509
rect 23112 28543 23164 28552
rect 23112 28509 23121 28543
rect 23121 28509 23155 28543
rect 23155 28509 23164 28543
rect 23112 28500 23164 28509
rect 23296 28543 23348 28552
rect 23296 28509 23305 28543
rect 23305 28509 23339 28543
rect 23339 28509 23348 28543
rect 32036 28568 32088 28620
rect 33692 28611 33744 28620
rect 33692 28577 33701 28611
rect 33701 28577 33735 28611
rect 33735 28577 33744 28611
rect 33692 28568 33744 28577
rect 34612 28568 34664 28620
rect 26884 28543 26936 28552
rect 23296 28500 23348 28509
rect 26884 28509 26893 28543
rect 26893 28509 26927 28543
rect 26927 28509 26936 28543
rect 26884 28500 26936 28509
rect 27068 28500 27120 28552
rect 27252 28500 27304 28552
rect 33416 28543 33468 28552
rect 18788 28432 18840 28484
rect 24768 28432 24820 28484
rect 33416 28509 33425 28543
rect 33425 28509 33459 28543
rect 33459 28509 33468 28543
rect 33416 28500 33468 28509
rect 33784 28543 33836 28552
rect 28172 28432 28224 28484
rect 28448 28432 28500 28484
rect 28816 28432 28868 28484
rect 33784 28509 33793 28543
rect 33793 28509 33827 28543
rect 33827 28509 33836 28543
rect 33784 28500 33836 28509
rect 33968 28543 34020 28552
rect 33968 28509 33977 28543
rect 33977 28509 34011 28543
rect 34011 28509 34020 28543
rect 33968 28500 34020 28509
rect 35808 28611 35860 28620
rect 35808 28577 35817 28611
rect 35817 28577 35851 28611
rect 35851 28577 35860 28611
rect 35808 28568 35860 28577
rect 37096 28611 37148 28620
rect 37096 28577 37105 28611
rect 37105 28577 37139 28611
rect 37139 28577 37148 28611
rect 37096 28568 37148 28577
rect 34796 28500 34848 28552
rect 38108 28543 38160 28552
rect 38108 28509 38117 28543
rect 38117 28509 38151 28543
rect 38151 28509 38160 28543
rect 38108 28500 38160 28509
rect 34520 28432 34572 28484
rect 16672 28364 16724 28416
rect 17592 28364 17644 28416
rect 32864 28364 32916 28416
rect 33416 28364 33468 28416
rect 36084 28364 36136 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 17316 28203 17368 28212
rect 17316 28169 17325 28203
rect 17325 28169 17359 28203
rect 17359 28169 17368 28203
rect 17316 28160 17368 28169
rect 23112 28160 23164 28212
rect 24768 28203 24820 28212
rect 24768 28169 24777 28203
rect 24777 28169 24811 28203
rect 24811 28169 24820 28203
rect 24768 28160 24820 28169
rect 27252 28203 27304 28212
rect 14188 28092 14240 28144
rect 20260 28092 20312 28144
rect 20628 28092 20680 28144
rect 21272 28092 21324 28144
rect 21916 28092 21968 28144
rect 12900 28067 12952 28076
rect 12900 28033 12909 28067
rect 12909 28033 12943 28067
rect 12943 28033 12952 28067
rect 12900 28024 12952 28033
rect 15292 28024 15344 28076
rect 17592 28067 17644 28076
rect 17592 28033 17601 28067
rect 17601 28033 17635 28067
rect 17635 28033 17644 28067
rect 17592 28024 17644 28033
rect 14464 27999 14516 28008
rect 14464 27965 14473 27999
rect 14473 27965 14507 27999
rect 14507 27965 14516 27999
rect 14464 27956 14516 27965
rect 15936 27999 15988 28008
rect 15936 27965 15945 27999
rect 15945 27965 15979 27999
rect 15979 27965 15988 27999
rect 15936 27956 15988 27965
rect 17776 28067 17828 28076
rect 17776 28033 17790 28067
rect 17790 28033 17824 28067
rect 17824 28033 17828 28067
rect 17776 28024 17828 28033
rect 18696 28024 18748 28076
rect 19432 28024 19484 28076
rect 20168 28067 20220 28076
rect 20168 28033 20202 28067
rect 20202 28033 20220 28067
rect 20168 28024 20220 28033
rect 20904 28024 20956 28076
rect 22284 28024 22336 28076
rect 27252 28169 27261 28203
rect 27261 28169 27295 28203
rect 27295 28169 27304 28203
rect 27252 28160 27304 28169
rect 28264 28203 28316 28212
rect 28264 28169 28273 28203
rect 28273 28169 28307 28203
rect 28307 28169 28316 28203
rect 28264 28160 28316 28169
rect 31760 28160 31812 28212
rect 33968 28160 34020 28212
rect 25320 28092 25372 28144
rect 25504 28092 25556 28144
rect 28448 28135 28500 28144
rect 28448 28101 28457 28135
rect 28457 28101 28491 28135
rect 28491 28101 28500 28135
rect 28448 28092 28500 28101
rect 22192 27956 22244 28008
rect 24308 27956 24360 28008
rect 17684 27888 17736 27940
rect 19432 27931 19484 27940
rect 19432 27897 19441 27931
rect 19441 27897 19475 27931
rect 19475 27897 19484 27931
rect 19432 27888 19484 27897
rect 25136 27956 25188 28008
rect 26884 28024 26936 28076
rect 27068 28067 27120 28076
rect 27068 28033 27077 28067
rect 27077 28033 27111 28067
rect 27111 28033 27120 28067
rect 28172 28067 28224 28076
rect 27068 28024 27120 28033
rect 28172 28033 28181 28067
rect 28181 28033 28215 28067
rect 28215 28033 28224 28067
rect 28172 28024 28224 28033
rect 28908 28067 28960 28076
rect 28908 28033 28917 28067
rect 28917 28033 28951 28067
rect 28951 28033 28960 28067
rect 28908 28024 28960 28033
rect 30380 28024 30432 28076
rect 31300 28067 31352 28076
rect 31300 28033 31309 28067
rect 31309 28033 31343 28067
rect 31343 28033 31352 28067
rect 31300 28024 31352 28033
rect 32956 28067 33008 28076
rect 32956 28033 32965 28067
rect 32965 28033 32999 28067
rect 32999 28033 33008 28067
rect 32956 28024 33008 28033
rect 33416 28024 33468 28076
rect 33784 28067 33836 28076
rect 33784 28033 33793 28067
rect 33793 28033 33827 28067
rect 33827 28033 33836 28067
rect 33784 28024 33836 28033
rect 34520 28024 34572 28076
rect 36728 28067 36780 28076
rect 36728 28033 36737 28067
rect 36737 28033 36771 28067
rect 36771 28033 36780 28067
rect 38384 28092 38436 28144
rect 36728 28024 36780 28033
rect 37556 28024 37608 28076
rect 27160 27956 27212 28008
rect 33692 27956 33744 28008
rect 31116 27888 31168 27940
rect 33508 27888 33560 27940
rect 35716 27999 35768 28008
rect 35716 27965 35725 27999
rect 35725 27965 35759 27999
rect 35759 27965 35768 27999
rect 35716 27956 35768 27965
rect 21272 27863 21324 27872
rect 21272 27829 21281 27863
rect 21281 27829 21315 27863
rect 21315 27829 21324 27863
rect 21272 27820 21324 27829
rect 22008 27863 22060 27872
rect 22008 27829 22017 27863
rect 22017 27829 22051 27863
rect 22051 27829 22060 27863
rect 22008 27820 22060 27829
rect 25412 27863 25464 27872
rect 25412 27829 25421 27863
rect 25421 27829 25455 27863
rect 25455 27829 25464 27863
rect 25412 27820 25464 27829
rect 29092 27863 29144 27872
rect 29092 27829 29101 27863
rect 29101 27829 29135 27863
rect 29135 27829 29144 27863
rect 29092 27820 29144 27829
rect 34060 27863 34112 27872
rect 34060 27829 34069 27863
rect 34069 27829 34103 27863
rect 34103 27829 34112 27863
rect 34060 27820 34112 27829
rect 37924 27820 37976 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 9588 27616 9640 27668
rect 14648 27616 14700 27668
rect 17776 27616 17828 27668
rect 20168 27659 20220 27668
rect 20168 27625 20177 27659
rect 20177 27625 20211 27659
rect 20211 27625 20220 27659
rect 20168 27616 20220 27625
rect 19432 27548 19484 27600
rect 22192 27616 22244 27668
rect 22284 27591 22336 27600
rect 22284 27557 22293 27591
rect 22293 27557 22327 27591
rect 22327 27557 22336 27591
rect 22284 27548 22336 27557
rect 27344 27591 27396 27600
rect 27344 27557 27353 27591
rect 27353 27557 27387 27591
rect 27387 27557 27396 27591
rect 27344 27548 27396 27557
rect 14832 27480 14884 27532
rect 17500 27480 17552 27532
rect 8392 27412 8444 27464
rect 12900 27412 12952 27464
rect 15292 27412 15344 27464
rect 17224 27412 17276 27464
rect 18420 27480 18472 27532
rect 20076 27480 20128 27532
rect 18328 27412 18380 27464
rect 19984 27412 20036 27464
rect 21272 27480 21324 27532
rect 22008 27523 22060 27532
rect 22008 27489 22017 27523
rect 22017 27489 22051 27523
rect 22051 27489 22060 27523
rect 22008 27480 22060 27489
rect 16764 27387 16816 27396
rect 16764 27353 16773 27387
rect 16773 27353 16807 27387
rect 16807 27353 16816 27387
rect 16764 27344 16816 27353
rect 17776 27344 17828 27396
rect 18788 27344 18840 27396
rect 20628 27455 20680 27464
rect 20628 27421 20637 27455
rect 20637 27421 20671 27455
rect 20671 27421 20680 27455
rect 20628 27412 20680 27421
rect 21456 27412 21508 27464
rect 22100 27412 22152 27464
rect 23204 27412 23256 27464
rect 26148 27412 26200 27464
rect 30840 27548 30892 27600
rect 32956 27548 33008 27600
rect 27712 27412 27764 27464
rect 28172 27412 28224 27464
rect 23020 27344 23072 27396
rect 27804 27344 27856 27396
rect 28264 27344 28316 27396
rect 7840 27319 7892 27328
rect 7840 27285 7849 27319
rect 7849 27285 7883 27319
rect 7883 27285 7892 27319
rect 7840 27276 7892 27285
rect 30748 27412 30800 27464
rect 33416 27480 33468 27532
rect 33508 27455 33560 27464
rect 30656 27276 30708 27328
rect 31392 27344 31444 27396
rect 33508 27421 33517 27455
rect 33517 27421 33551 27455
rect 33551 27421 33560 27455
rect 33508 27412 33560 27421
rect 37188 27523 37240 27532
rect 37188 27489 37197 27523
rect 37197 27489 37231 27523
rect 37231 27489 37240 27523
rect 37188 27480 37240 27489
rect 37924 27523 37976 27532
rect 37924 27489 37933 27523
rect 37933 27489 37967 27523
rect 37967 27489 37976 27523
rect 37924 27480 37976 27489
rect 38108 27523 38160 27532
rect 38108 27489 38117 27523
rect 38117 27489 38151 27523
rect 38151 27489 38160 27523
rect 38108 27480 38160 27489
rect 33324 27319 33376 27328
rect 33324 27285 33333 27319
rect 33333 27285 33367 27319
rect 33367 27285 33376 27319
rect 33324 27276 33376 27285
rect 34796 27344 34848 27396
rect 37556 27276 37608 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 8024 27072 8076 27124
rect 17224 27115 17276 27124
rect 17224 27081 17233 27115
rect 17233 27081 17267 27115
rect 17267 27081 17276 27115
rect 17224 27072 17276 27081
rect 17776 27115 17828 27124
rect 17776 27081 17785 27115
rect 17785 27081 17819 27115
rect 17819 27081 17828 27115
rect 17776 27072 17828 27081
rect 18512 27115 18564 27124
rect 18512 27081 18521 27115
rect 18521 27081 18555 27115
rect 18555 27081 18564 27115
rect 18512 27072 18564 27081
rect 20260 27047 20312 27056
rect 20260 27013 20269 27047
rect 20269 27013 20303 27047
rect 20303 27013 20312 27047
rect 20260 27004 20312 27013
rect 22376 27004 22428 27056
rect 26240 27004 26292 27056
rect 29092 27004 29144 27056
rect 7840 26936 7892 26988
rect 14924 26979 14976 26988
rect 14924 26945 14933 26979
rect 14933 26945 14967 26979
rect 14967 26945 14976 26979
rect 14924 26936 14976 26945
rect 16856 26979 16908 26988
rect 16856 26945 16865 26979
rect 16865 26945 16899 26979
rect 16899 26945 16908 26979
rect 16856 26936 16908 26945
rect 15476 26911 15528 26920
rect 15476 26877 15485 26911
rect 15485 26877 15519 26911
rect 15519 26877 15528 26911
rect 15476 26868 15528 26877
rect 18052 26868 18104 26920
rect 20076 26936 20128 26988
rect 21824 26979 21876 26988
rect 21824 26945 21833 26979
rect 21833 26945 21867 26979
rect 21867 26945 21876 26979
rect 21824 26936 21876 26945
rect 18788 26911 18840 26920
rect 18788 26877 18797 26911
rect 18797 26877 18831 26911
rect 18831 26877 18840 26911
rect 22008 26936 22060 26988
rect 22284 26936 22336 26988
rect 23204 26979 23256 26988
rect 23204 26945 23213 26979
rect 23213 26945 23247 26979
rect 23247 26945 23256 26979
rect 23204 26936 23256 26945
rect 25412 26979 25464 26988
rect 18788 26868 18840 26877
rect 23388 26868 23440 26920
rect 20168 26800 20220 26852
rect 22100 26800 22152 26852
rect 25412 26945 25421 26979
rect 25421 26945 25455 26979
rect 25455 26945 25464 26979
rect 25412 26936 25464 26945
rect 25872 26979 25924 26988
rect 25872 26945 25881 26979
rect 25881 26945 25915 26979
rect 25915 26945 25924 26979
rect 25872 26936 25924 26945
rect 26148 26979 26200 26988
rect 26148 26945 26157 26979
rect 26157 26945 26191 26979
rect 26191 26945 26200 26979
rect 26148 26936 26200 26945
rect 27344 26979 27396 26988
rect 27344 26945 27353 26979
rect 27353 26945 27387 26979
rect 27387 26945 27396 26979
rect 27344 26936 27396 26945
rect 27712 26936 27764 26988
rect 35716 27004 35768 27056
rect 30380 26979 30432 26988
rect 26056 26868 26108 26920
rect 27620 26911 27672 26920
rect 27620 26877 27629 26911
rect 27629 26877 27663 26911
rect 27663 26877 27672 26911
rect 27620 26868 27672 26877
rect 26700 26800 26752 26852
rect 30380 26945 30389 26979
rect 30389 26945 30423 26979
rect 30423 26945 30432 26979
rect 30380 26936 30432 26945
rect 30564 26979 30616 26988
rect 30564 26945 30573 26979
rect 30573 26945 30607 26979
rect 30607 26945 30616 26979
rect 30564 26936 30616 26945
rect 30840 26936 30892 26988
rect 34152 26936 34204 26988
rect 36176 27004 36228 27056
rect 37372 26936 37424 26988
rect 29828 26911 29880 26920
rect 29828 26877 29837 26911
rect 29837 26877 29871 26911
rect 29871 26877 29880 26911
rect 29828 26868 29880 26877
rect 30656 26868 30708 26920
rect 30932 26868 30984 26920
rect 37464 26868 37516 26920
rect 37740 26868 37792 26920
rect 28448 26843 28500 26852
rect 28448 26809 28457 26843
rect 28457 26809 28491 26843
rect 28491 26809 28500 26843
rect 28448 26800 28500 26809
rect 21180 26775 21232 26784
rect 21180 26741 21189 26775
rect 21189 26741 21223 26775
rect 21223 26741 21232 26775
rect 21180 26732 21232 26741
rect 22008 26732 22060 26784
rect 22928 26732 22980 26784
rect 24952 26775 25004 26784
rect 24952 26741 24961 26775
rect 24961 26741 24995 26775
rect 24995 26741 25004 26775
rect 24952 26732 25004 26741
rect 25320 26775 25372 26784
rect 25320 26741 25329 26775
rect 25329 26741 25363 26775
rect 25363 26741 25372 26775
rect 25320 26732 25372 26741
rect 25872 26732 25924 26784
rect 27160 26775 27212 26784
rect 27160 26741 27169 26775
rect 27169 26741 27203 26775
rect 27203 26741 27212 26775
rect 27160 26732 27212 26741
rect 32036 26732 32088 26784
rect 32772 26732 32824 26784
rect 33508 26732 33560 26784
rect 34520 26732 34572 26784
rect 35624 26732 35676 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 15200 26528 15252 26580
rect 15476 26528 15528 26580
rect 16856 26460 16908 26512
rect 18788 26528 18840 26580
rect 20628 26528 20680 26580
rect 26056 26571 26108 26580
rect 16580 26392 16632 26444
rect 16212 26324 16264 26376
rect 17040 26367 17092 26376
rect 17040 26333 17049 26367
rect 17049 26333 17083 26367
rect 17083 26333 17092 26367
rect 17040 26324 17092 26333
rect 23388 26460 23440 26512
rect 26056 26537 26065 26571
rect 26065 26537 26099 26571
rect 26099 26537 26108 26571
rect 26056 26528 26108 26537
rect 27804 26528 27856 26580
rect 31392 26571 31444 26580
rect 31392 26537 31401 26571
rect 31401 26537 31435 26571
rect 31435 26537 31444 26571
rect 31392 26528 31444 26537
rect 26700 26460 26752 26512
rect 30656 26460 30708 26512
rect 32956 26528 33008 26580
rect 34152 26571 34204 26580
rect 34152 26537 34161 26571
rect 34161 26537 34195 26571
rect 34195 26537 34204 26571
rect 34152 26528 34204 26537
rect 19340 26392 19392 26444
rect 20076 26392 20128 26444
rect 20260 26392 20312 26444
rect 18052 26324 18104 26376
rect 18328 26367 18380 26376
rect 18328 26333 18337 26367
rect 18337 26333 18371 26367
rect 18371 26333 18380 26367
rect 18328 26324 18380 26333
rect 16856 26299 16908 26308
rect 16856 26265 16865 26299
rect 16865 26265 16899 26299
rect 16899 26265 16908 26299
rect 16856 26256 16908 26265
rect 18512 26299 18564 26308
rect 18512 26265 18521 26299
rect 18521 26265 18555 26299
rect 18555 26265 18564 26299
rect 18512 26256 18564 26265
rect 19248 26299 19300 26308
rect 19248 26265 19257 26299
rect 19257 26265 19291 26299
rect 19291 26265 19300 26299
rect 19248 26256 19300 26265
rect 16948 26188 17000 26240
rect 21088 26324 21140 26376
rect 21180 26324 21232 26376
rect 23480 26324 23532 26376
rect 24400 26324 24452 26376
rect 24952 26367 25004 26376
rect 24952 26333 24986 26367
rect 24986 26333 25004 26367
rect 24952 26324 25004 26333
rect 29828 26324 29880 26376
rect 30564 26367 30616 26376
rect 30564 26333 30573 26367
rect 30573 26333 30607 26367
rect 30607 26333 30616 26367
rect 30564 26324 30616 26333
rect 31668 26367 31720 26376
rect 31668 26333 31677 26367
rect 31677 26333 31711 26367
rect 31711 26333 31720 26367
rect 31668 26324 31720 26333
rect 32128 26392 32180 26444
rect 32036 26367 32088 26376
rect 20812 26256 20864 26308
rect 21824 26256 21876 26308
rect 22744 26256 22796 26308
rect 27160 26256 27212 26308
rect 32036 26333 32045 26367
rect 32045 26333 32079 26367
rect 32079 26333 32088 26367
rect 32036 26324 32088 26333
rect 33324 26392 33376 26444
rect 32864 26367 32916 26376
rect 32864 26333 32873 26367
rect 32873 26333 32907 26367
rect 32907 26333 32916 26367
rect 32864 26324 32916 26333
rect 33048 26324 33100 26376
rect 33508 26367 33560 26376
rect 33508 26333 33517 26367
rect 33517 26333 33551 26367
rect 33551 26333 33560 26367
rect 34520 26392 34572 26444
rect 34704 26392 34756 26444
rect 35348 26392 35400 26444
rect 36084 26435 36136 26444
rect 36084 26401 36093 26435
rect 36093 26401 36127 26435
rect 36127 26401 36136 26435
rect 36084 26392 36136 26401
rect 33508 26324 33560 26333
rect 33232 26256 33284 26308
rect 34060 26324 34112 26376
rect 34980 26367 35032 26376
rect 34980 26333 34989 26367
rect 34989 26333 35023 26367
rect 35023 26333 35032 26367
rect 36176 26367 36228 26376
rect 34980 26324 35032 26333
rect 36176 26333 36185 26367
rect 36185 26333 36219 26367
rect 36219 26333 36228 26367
rect 36176 26324 36228 26333
rect 37372 26367 37424 26376
rect 37372 26333 37381 26367
rect 37381 26333 37415 26367
rect 37415 26333 37424 26367
rect 37372 26324 37424 26333
rect 37464 26299 37516 26308
rect 37464 26265 37473 26299
rect 37473 26265 37507 26299
rect 37507 26265 37516 26299
rect 37464 26256 37516 26265
rect 22008 26188 22060 26240
rect 30472 26188 30524 26240
rect 31484 26188 31536 26240
rect 34520 26188 34572 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 17040 26027 17092 26036
rect 17040 25993 17049 26027
rect 17049 25993 17083 26027
rect 17083 25993 17092 26027
rect 17040 25984 17092 25993
rect 18328 25984 18380 26036
rect 20904 25984 20956 26036
rect 21088 25984 21140 26036
rect 21272 25984 21324 26036
rect 22744 26027 22796 26036
rect 22744 25993 22753 26027
rect 22753 25993 22787 26027
rect 22787 25993 22796 26027
rect 22744 25984 22796 25993
rect 15844 25916 15896 25968
rect 31852 25984 31904 26036
rect 32128 25984 32180 26036
rect 33048 25984 33100 26036
rect 33232 26027 33284 26036
rect 33232 25993 33241 26027
rect 33241 25993 33275 26027
rect 33275 25993 33284 26027
rect 33232 25984 33284 25993
rect 34980 25984 35032 26036
rect 16672 25891 16724 25900
rect 16672 25857 16681 25891
rect 16681 25857 16715 25891
rect 16715 25857 16724 25891
rect 16672 25848 16724 25857
rect 16948 25848 17000 25900
rect 19156 25848 19208 25900
rect 20904 25891 20956 25900
rect 16580 25780 16632 25832
rect 17868 25780 17920 25832
rect 19432 25780 19484 25832
rect 20904 25857 20913 25891
rect 20913 25857 20947 25891
rect 20947 25857 20956 25891
rect 20904 25848 20956 25857
rect 21824 25891 21876 25900
rect 21824 25857 21833 25891
rect 21833 25857 21867 25891
rect 21867 25857 21876 25891
rect 21824 25848 21876 25857
rect 22008 25891 22060 25900
rect 22008 25857 22017 25891
rect 22017 25857 22051 25891
rect 22051 25857 22060 25891
rect 22008 25848 22060 25857
rect 22928 25891 22980 25900
rect 22928 25857 22937 25891
rect 22937 25857 22971 25891
rect 22971 25857 22980 25891
rect 22928 25848 22980 25857
rect 23020 25848 23072 25900
rect 25044 25891 25096 25900
rect 25044 25857 25053 25891
rect 25053 25857 25087 25891
rect 25087 25857 25096 25891
rect 25044 25848 25096 25857
rect 30656 25848 30708 25900
rect 31852 25848 31904 25900
rect 20812 25780 20864 25832
rect 23388 25780 23440 25832
rect 25320 25823 25372 25832
rect 25320 25789 25329 25823
rect 25329 25789 25363 25823
rect 25363 25789 25372 25823
rect 25320 25780 25372 25789
rect 30932 25780 30984 25832
rect 31484 25823 31536 25832
rect 31484 25789 31493 25823
rect 31493 25789 31527 25823
rect 31527 25789 31536 25823
rect 32220 25823 32272 25832
rect 31484 25780 31536 25789
rect 32220 25789 32229 25823
rect 32229 25789 32263 25823
rect 32263 25789 32272 25823
rect 32220 25780 32272 25789
rect 22836 25712 22888 25764
rect 23112 25712 23164 25764
rect 33784 25848 33836 25900
rect 34520 25891 34572 25900
rect 34520 25857 34529 25891
rect 34529 25857 34563 25891
rect 34563 25857 34572 25891
rect 34520 25848 34572 25857
rect 34796 25848 34848 25900
rect 34980 25848 35032 25900
rect 35348 25891 35400 25900
rect 35348 25857 35357 25891
rect 35357 25857 35391 25891
rect 35391 25857 35400 25891
rect 35348 25848 35400 25857
rect 16212 25644 16264 25696
rect 19064 25687 19116 25696
rect 19064 25653 19073 25687
rect 19073 25653 19107 25687
rect 19107 25653 19116 25687
rect 19064 25644 19116 25653
rect 19340 25644 19392 25696
rect 29184 25687 29236 25696
rect 29184 25653 29193 25687
rect 29193 25653 29227 25687
rect 29227 25653 29236 25687
rect 29184 25644 29236 25653
rect 34704 25644 34756 25696
rect 36544 25687 36596 25696
rect 36544 25653 36553 25687
rect 36553 25653 36587 25687
rect 36587 25653 36596 25687
rect 36544 25644 36596 25653
rect 37924 25644 37976 25696
rect 38108 25687 38160 25696
rect 38108 25653 38117 25687
rect 38117 25653 38151 25687
rect 38151 25653 38160 25687
rect 38108 25644 38160 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 18052 25483 18104 25492
rect 18052 25449 18061 25483
rect 18061 25449 18095 25483
rect 18095 25449 18104 25483
rect 18052 25440 18104 25449
rect 18512 25440 18564 25492
rect 25044 25440 25096 25492
rect 32220 25483 32272 25492
rect 32220 25449 32229 25483
rect 32229 25449 32263 25483
rect 32263 25449 32272 25483
rect 32220 25440 32272 25449
rect 16948 25372 17000 25424
rect 18328 25347 18380 25356
rect 18328 25313 18337 25347
rect 18337 25313 18371 25347
rect 18371 25313 18380 25347
rect 18328 25304 18380 25313
rect 19984 25372 20036 25424
rect 34520 25372 34572 25424
rect 19064 25304 19116 25356
rect 22008 25304 22060 25356
rect 24400 25347 24452 25356
rect 24400 25313 24409 25347
rect 24409 25313 24443 25347
rect 24443 25313 24452 25347
rect 24400 25304 24452 25313
rect 34796 25304 34848 25356
rect 37188 25347 37240 25356
rect 37188 25313 37197 25347
rect 37197 25313 37231 25347
rect 37231 25313 37240 25347
rect 37188 25304 37240 25313
rect 37924 25347 37976 25356
rect 37924 25313 37933 25347
rect 37933 25313 37967 25347
rect 37967 25313 37976 25347
rect 37924 25304 37976 25313
rect 38108 25347 38160 25356
rect 38108 25313 38117 25347
rect 38117 25313 38151 25347
rect 38151 25313 38160 25347
rect 38108 25304 38160 25313
rect 16580 25279 16632 25288
rect 16580 25245 16589 25279
rect 16589 25245 16623 25279
rect 16623 25245 16632 25279
rect 16580 25236 16632 25245
rect 18236 25279 18288 25288
rect 18236 25245 18245 25279
rect 18245 25245 18279 25279
rect 18279 25245 18288 25279
rect 18236 25236 18288 25245
rect 19340 25236 19392 25288
rect 20720 25279 20772 25288
rect 20720 25245 20729 25279
rect 20729 25245 20763 25279
rect 20763 25245 20772 25279
rect 20720 25236 20772 25245
rect 20812 25279 20864 25288
rect 20812 25245 20821 25279
rect 20821 25245 20855 25279
rect 20855 25245 20864 25279
rect 20812 25236 20864 25245
rect 20996 25279 21048 25288
rect 20996 25245 21005 25279
rect 21005 25245 21039 25279
rect 21039 25245 21048 25279
rect 20996 25236 21048 25245
rect 29184 25236 29236 25288
rect 29828 25236 29880 25288
rect 32036 25279 32088 25288
rect 32036 25245 32045 25279
rect 32045 25245 32079 25279
rect 32079 25245 32088 25279
rect 32036 25236 32088 25245
rect 32864 25236 32916 25288
rect 34888 25279 34940 25288
rect 34888 25245 34897 25279
rect 34897 25245 34931 25279
rect 34931 25245 34940 25279
rect 34888 25236 34940 25245
rect 35348 25236 35400 25288
rect 24492 25168 24544 25220
rect 19156 25100 19208 25152
rect 30472 25143 30524 25152
rect 30472 25109 30481 25143
rect 30481 25109 30515 25143
rect 30515 25109 30524 25143
rect 30472 25100 30524 25109
rect 34796 25100 34848 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 15660 24803 15712 24812
rect 15660 24769 15669 24803
rect 15669 24769 15703 24803
rect 15703 24769 15712 24803
rect 15660 24760 15712 24769
rect 16856 24760 16908 24812
rect 17868 24760 17920 24812
rect 20720 24760 20772 24812
rect 24492 24939 24544 24948
rect 24492 24905 24501 24939
rect 24501 24905 24535 24939
rect 24535 24905 24544 24939
rect 24492 24896 24544 24905
rect 32036 24896 32088 24948
rect 21088 24760 21140 24812
rect 34888 24896 34940 24948
rect 21272 24803 21324 24812
rect 21272 24769 21281 24803
rect 21281 24769 21315 24803
rect 21315 24769 21324 24803
rect 21272 24760 21324 24769
rect 20536 24692 20588 24744
rect 21640 24692 21692 24744
rect 25320 24760 25372 24812
rect 27344 24760 27396 24812
rect 25688 24692 25740 24744
rect 27988 24760 28040 24812
rect 31760 24760 31812 24812
rect 30012 24692 30064 24744
rect 32956 24760 33008 24812
rect 33968 24692 34020 24744
rect 34152 24803 34204 24812
rect 34152 24769 34161 24803
rect 34161 24769 34195 24803
rect 34195 24769 34204 24803
rect 34152 24760 34204 24769
rect 34520 24692 34572 24744
rect 35900 24803 35952 24812
rect 35900 24769 35909 24803
rect 35909 24769 35943 24803
rect 35943 24769 35952 24803
rect 35900 24760 35952 24769
rect 36084 24692 36136 24744
rect 29092 24624 29144 24676
rect 33600 24624 33652 24676
rect 15936 24556 15988 24608
rect 20444 24556 20496 24608
rect 21272 24556 21324 24608
rect 22192 24599 22244 24608
rect 22192 24565 22201 24599
rect 22201 24565 22235 24599
rect 22235 24565 22244 24599
rect 22192 24556 22244 24565
rect 28080 24599 28132 24608
rect 28080 24565 28089 24599
rect 28089 24565 28123 24599
rect 28123 24565 28132 24599
rect 28080 24556 28132 24565
rect 29736 24556 29788 24608
rect 30472 24556 30524 24608
rect 33692 24556 33744 24608
rect 34152 24556 34204 24608
rect 34704 24556 34756 24608
rect 37832 24599 37884 24608
rect 37832 24565 37841 24599
rect 37841 24565 37875 24599
rect 37875 24565 37884 24599
rect 37832 24556 37884 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 15660 24352 15712 24404
rect 15476 24191 15528 24200
rect 15476 24157 15485 24191
rect 15485 24157 15519 24191
rect 15519 24157 15528 24191
rect 15476 24148 15528 24157
rect 20996 24352 21048 24404
rect 21180 24352 21232 24404
rect 19248 24216 19300 24268
rect 16856 24148 16908 24200
rect 18236 24191 18288 24200
rect 18236 24157 18245 24191
rect 18245 24157 18279 24191
rect 18279 24157 18288 24191
rect 18236 24148 18288 24157
rect 20168 24148 20220 24200
rect 20444 24191 20496 24200
rect 20444 24157 20453 24191
rect 20453 24157 20487 24191
rect 20487 24157 20496 24191
rect 20444 24148 20496 24157
rect 21640 24216 21692 24268
rect 16948 24080 17000 24132
rect 16028 24012 16080 24064
rect 18328 24012 18380 24064
rect 33140 24352 33192 24404
rect 33416 24352 33468 24404
rect 35348 24352 35400 24404
rect 35624 24395 35676 24404
rect 35624 24361 35633 24395
rect 35633 24361 35667 24395
rect 35667 24361 35676 24395
rect 35624 24352 35676 24361
rect 22192 24284 22244 24336
rect 27344 24327 27396 24336
rect 27344 24293 27353 24327
rect 27353 24293 27387 24327
rect 27387 24293 27396 24327
rect 27344 24284 27396 24293
rect 22284 24259 22336 24268
rect 22284 24225 22293 24259
rect 22293 24225 22327 24259
rect 22327 24225 22336 24259
rect 22284 24216 22336 24225
rect 25688 24259 25740 24268
rect 25688 24225 25697 24259
rect 25697 24225 25731 24259
rect 25731 24225 25740 24259
rect 25688 24216 25740 24225
rect 31760 24216 31812 24268
rect 33692 24259 33744 24268
rect 33692 24225 33701 24259
rect 33701 24225 33735 24259
rect 33735 24225 33744 24259
rect 33692 24216 33744 24225
rect 33784 24259 33836 24268
rect 33784 24225 33793 24259
rect 33793 24225 33827 24259
rect 33827 24225 33836 24259
rect 33784 24216 33836 24225
rect 36084 24216 36136 24268
rect 36544 24216 36596 24268
rect 38108 24259 38160 24268
rect 38108 24225 38117 24259
rect 38117 24225 38151 24259
rect 38151 24225 38160 24259
rect 38108 24216 38160 24225
rect 22008 24012 22060 24064
rect 26792 24148 26844 24200
rect 26976 24148 27028 24200
rect 28080 24148 28132 24200
rect 29552 24191 29604 24200
rect 26608 24123 26660 24132
rect 26608 24089 26617 24123
rect 26617 24089 26651 24123
rect 26651 24089 26660 24123
rect 26608 24080 26660 24089
rect 28540 24080 28592 24132
rect 29552 24157 29561 24191
rect 29561 24157 29595 24191
rect 29595 24157 29604 24191
rect 29552 24148 29604 24157
rect 29736 24191 29788 24200
rect 29736 24157 29743 24191
rect 29743 24157 29788 24191
rect 29736 24148 29788 24157
rect 29920 24191 29972 24200
rect 29920 24157 29929 24191
rect 29929 24157 29963 24191
rect 29963 24157 29972 24191
rect 29920 24148 29972 24157
rect 30012 24191 30064 24200
rect 30012 24157 30026 24191
rect 30026 24157 30060 24191
rect 30060 24157 30064 24191
rect 30012 24148 30064 24157
rect 30748 24148 30800 24200
rect 33416 24191 33468 24200
rect 33416 24157 33425 24191
rect 33425 24157 33459 24191
rect 33459 24157 33468 24191
rect 33416 24148 33468 24157
rect 33600 24191 33652 24200
rect 33600 24157 33609 24191
rect 33609 24157 33643 24191
rect 33643 24157 33652 24191
rect 33600 24148 33652 24157
rect 35440 24191 35492 24200
rect 30104 24080 30156 24132
rect 31024 24080 31076 24132
rect 35440 24157 35449 24191
rect 35449 24157 35483 24191
rect 35483 24157 35492 24191
rect 35440 24148 35492 24157
rect 35900 24148 35952 24200
rect 37464 24080 37516 24132
rect 22652 24055 22704 24064
rect 22652 24021 22661 24055
rect 22661 24021 22695 24055
rect 22695 24021 22704 24055
rect 22652 24012 22704 24021
rect 25964 24055 26016 24064
rect 25964 24021 25973 24055
rect 25973 24021 26007 24055
rect 26007 24021 26016 24055
rect 25964 24012 26016 24021
rect 27344 24012 27396 24064
rect 30196 24055 30248 24064
rect 30196 24021 30205 24055
rect 30205 24021 30239 24055
rect 30239 24021 30248 24055
rect 30196 24012 30248 24021
rect 30748 24055 30800 24064
rect 30748 24021 30757 24055
rect 30757 24021 30791 24055
rect 30791 24021 30800 24055
rect 30748 24012 30800 24021
rect 32680 24012 32732 24064
rect 35532 24012 35584 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 15936 23851 15988 23860
rect 15936 23817 15945 23851
rect 15945 23817 15979 23851
rect 15979 23817 15988 23851
rect 15936 23808 15988 23817
rect 18236 23808 18288 23860
rect 18420 23851 18472 23860
rect 18420 23817 18429 23851
rect 18429 23817 18463 23851
rect 18463 23817 18472 23851
rect 18420 23808 18472 23817
rect 21088 23851 21140 23860
rect 21088 23817 21097 23851
rect 21097 23817 21131 23851
rect 21131 23817 21140 23851
rect 21088 23808 21140 23817
rect 22008 23808 22060 23860
rect 27344 23808 27396 23860
rect 27988 23808 28040 23860
rect 28540 23808 28592 23860
rect 30748 23808 30800 23860
rect 16304 23740 16356 23792
rect 18328 23783 18380 23792
rect 15844 23672 15896 23724
rect 16028 23715 16080 23724
rect 16028 23681 16037 23715
rect 16037 23681 16071 23715
rect 16071 23681 16080 23715
rect 16028 23672 16080 23681
rect 17500 23672 17552 23724
rect 18328 23749 18337 23783
rect 18337 23749 18371 23783
rect 18371 23749 18380 23783
rect 18328 23740 18380 23749
rect 20168 23740 20220 23792
rect 22652 23740 22704 23792
rect 25964 23740 26016 23792
rect 17868 23604 17920 23656
rect 19432 23715 19484 23724
rect 19432 23681 19441 23715
rect 19441 23681 19475 23715
rect 19475 23681 19484 23715
rect 19432 23672 19484 23681
rect 20904 23715 20956 23724
rect 20904 23681 20913 23715
rect 20913 23681 20947 23715
rect 20947 23681 20956 23715
rect 20904 23672 20956 23681
rect 21180 23672 21232 23724
rect 22100 23672 22152 23724
rect 24308 23672 24360 23724
rect 26976 23715 27028 23724
rect 26976 23681 26985 23715
rect 26985 23681 27019 23715
rect 27019 23681 27028 23715
rect 26976 23672 27028 23681
rect 27896 23715 27948 23724
rect 27896 23681 27905 23715
rect 27905 23681 27939 23715
rect 27939 23681 27948 23715
rect 27896 23672 27948 23681
rect 25044 23647 25096 23656
rect 25044 23613 25053 23647
rect 25053 23613 25087 23647
rect 25087 23613 25096 23647
rect 25044 23604 25096 23613
rect 26608 23604 26660 23656
rect 27436 23604 27488 23656
rect 29000 23672 29052 23724
rect 32312 23740 32364 23792
rect 32956 23740 33008 23792
rect 34520 23808 34572 23860
rect 35624 23808 35676 23860
rect 35900 23808 35952 23860
rect 35532 23783 35584 23792
rect 29920 23715 29972 23724
rect 29920 23681 29929 23715
rect 29929 23681 29963 23715
rect 29963 23681 29972 23715
rect 29920 23672 29972 23681
rect 30012 23715 30064 23724
rect 30012 23681 30021 23715
rect 30021 23681 30055 23715
rect 30055 23681 30064 23715
rect 30196 23715 30248 23724
rect 30012 23672 30064 23681
rect 30196 23681 30205 23715
rect 30205 23681 30239 23715
rect 30239 23681 30248 23715
rect 30196 23672 30248 23681
rect 33600 23715 33652 23724
rect 33600 23681 33609 23715
rect 33609 23681 33643 23715
rect 33643 23681 33652 23715
rect 33600 23672 33652 23681
rect 34060 23672 34112 23724
rect 35532 23749 35566 23783
rect 35566 23749 35584 23783
rect 35532 23740 35584 23749
rect 28816 23604 28868 23656
rect 33968 23604 34020 23656
rect 29092 23536 29144 23588
rect 30104 23536 30156 23588
rect 32864 23536 32916 23588
rect 15568 23511 15620 23520
rect 15568 23477 15577 23511
rect 15577 23477 15611 23511
rect 15611 23477 15620 23511
rect 15568 23468 15620 23477
rect 15660 23511 15712 23520
rect 15660 23477 15669 23511
rect 15669 23477 15703 23511
rect 15703 23477 15712 23511
rect 18696 23511 18748 23520
rect 15660 23468 15712 23477
rect 18696 23477 18705 23511
rect 18705 23477 18739 23511
rect 18739 23477 18748 23511
rect 18696 23468 18748 23477
rect 29644 23468 29696 23520
rect 32680 23468 32732 23520
rect 35348 23672 35400 23724
rect 37280 23672 37332 23724
rect 38292 23672 38344 23724
rect 37924 23468 37976 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 15660 23264 15712 23316
rect 17500 23264 17552 23316
rect 26792 23264 26844 23316
rect 27344 23264 27396 23316
rect 29552 23264 29604 23316
rect 15476 23196 15528 23248
rect 1768 23103 1820 23112
rect 1768 23069 1777 23103
rect 1777 23069 1811 23103
rect 1811 23069 1820 23103
rect 1768 23060 1820 23069
rect 14188 23060 14240 23112
rect 15568 23060 15620 23112
rect 16304 23103 16356 23112
rect 16304 23069 16313 23103
rect 16313 23069 16347 23103
rect 16347 23069 16356 23103
rect 16304 23060 16356 23069
rect 16488 23103 16540 23112
rect 16488 23069 16497 23103
rect 16497 23069 16531 23103
rect 16531 23069 16540 23103
rect 19432 23103 19484 23112
rect 16488 23060 16540 23069
rect 19432 23069 19441 23103
rect 19441 23069 19475 23103
rect 19475 23069 19484 23103
rect 19432 23060 19484 23069
rect 22008 23060 22060 23112
rect 22100 23103 22152 23112
rect 22100 23069 22109 23103
rect 22109 23069 22143 23103
rect 22143 23069 22152 23103
rect 22100 23060 22152 23069
rect 25044 23060 25096 23112
rect 28264 23060 28316 23112
rect 28816 23103 28868 23112
rect 28816 23069 28825 23103
rect 28825 23069 28859 23103
rect 28859 23069 28868 23103
rect 28816 23060 28868 23069
rect 29000 23103 29052 23112
rect 29000 23069 29009 23103
rect 29009 23069 29043 23103
rect 29043 23069 29052 23103
rect 29000 23060 29052 23069
rect 29828 23060 29880 23112
rect 30104 23196 30156 23248
rect 33784 23239 33836 23248
rect 33784 23205 33793 23239
rect 33793 23205 33827 23239
rect 33827 23205 33836 23239
rect 33784 23196 33836 23205
rect 37832 23196 37884 23248
rect 37188 23171 37240 23180
rect 37188 23137 37197 23171
rect 37197 23137 37231 23171
rect 37231 23137 37240 23171
rect 37188 23128 37240 23137
rect 37924 23171 37976 23180
rect 37924 23137 37933 23171
rect 37933 23137 37967 23171
rect 37967 23137 37976 23171
rect 37924 23128 37976 23137
rect 30104 23103 30156 23112
rect 30104 23069 30113 23103
rect 30113 23069 30147 23103
rect 30147 23069 30156 23103
rect 30104 23060 30156 23069
rect 30932 23060 30984 23112
rect 32680 23060 32732 23112
rect 33600 23103 33652 23112
rect 33600 23069 33609 23103
rect 33609 23069 33643 23103
rect 33643 23069 33652 23103
rect 33600 23060 33652 23069
rect 35440 23103 35492 23112
rect 35440 23069 35449 23103
rect 35449 23069 35483 23103
rect 35483 23069 35492 23103
rect 35440 23060 35492 23069
rect 9588 22992 9640 23044
rect 14556 22992 14608 23044
rect 24676 23035 24728 23044
rect 24676 23001 24710 23035
rect 24710 23001 24728 23035
rect 27436 23035 27488 23044
rect 24676 22992 24728 23001
rect 27436 23001 27445 23035
rect 27445 23001 27479 23035
rect 27479 23001 27488 23035
rect 27436 22992 27488 23001
rect 28908 22992 28960 23044
rect 1952 22924 2004 22976
rect 20904 22924 20956 22976
rect 21640 22924 21692 22976
rect 22008 22924 22060 22976
rect 25780 22967 25832 22976
rect 25780 22933 25789 22967
rect 25789 22933 25823 22967
rect 25823 22933 25832 22967
rect 25780 22924 25832 22933
rect 26976 22924 27028 22976
rect 29736 22924 29788 22976
rect 32128 22992 32180 23044
rect 31024 22924 31076 22976
rect 31208 22967 31260 22976
rect 31208 22933 31217 22967
rect 31217 22933 31251 22967
rect 31251 22933 31260 22967
rect 31208 22924 31260 22933
rect 35532 22924 35584 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 19432 22720 19484 22772
rect 20812 22720 20864 22772
rect 24676 22763 24728 22772
rect 24676 22729 24685 22763
rect 24685 22729 24719 22763
rect 24719 22729 24728 22763
rect 24676 22720 24728 22729
rect 32128 22763 32180 22772
rect 32128 22729 32137 22763
rect 32137 22729 32171 22763
rect 32171 22729 32180 22763
rect 32128 22720 32180 22729
rect 33600 22720 33652 22772
rect 1952 22695 2004 22704
rect 1952 22661 1961 22695
rect 1961 22661 1995 22695
rect 1995 22661 2004 22695
rect 1952 22652 2004 22661
rect 18696 22652 18748 22704
rect 22376 22695 22428 22704
rect 22376 22661 22385 22695
rect 22385 22661 22419 22695
rect 22419 22661 22428 22695
rect 22376 22652 22428 22661
rect 1768 22627 1820 22636
rect 1768 22593 1777 22627
rect 1777 22593 1811 22627
rect 1811 22593 1820 22627
rect 1768 22584 1820 22593
rect 16488 22584 16540 22636
rect 21640 22584 21692 22636
rect 23112 22627 23164 22636
rect 23112 22593 23121 22627
rect 23121 22593 23155 22627
rect 23155 22593 23164 22627
rect 23112 22584 23164 22593
rect 24952 22652 25004 22704
rect 25688 22652 25740 22704
rect 28908 22652 28960 22704
rect 2780 22559 2832 22568
rect 2780 22525 2789 22559
rect 2789 22525 2823 22559
rect 2823 22525 2832 22559
rect 2780 22516 2832 22525
rect 17868 22559 17920 22568
rect 17868 22525 17877 22559
rect 17877 22525 17911 22559
rect 17911 22525 17920 22559
rect 17868 22516 17920 22525
rect 20536 22559 20588 22568
rect 20536 22525 20545 22559
rect 20545 22525 20579 22559
rect 20579 22525 20588 22559
rect 20536 22516 20588 22525
rect 23296 22516 23348 22568
rect 25780 22584 25832 22636
rect 28264 22584 28316 22636
rect 29644 22627 29696 22636
rect 29644 22593 29653 22627
rect 29653 22593 29687 22627
rect 29687 22593 29696 22627
rect 29644 22584 29696 22593
rect 29736 22627 29788 22636
rect 29736 22593 29745 22627
rect 29745 22593 29779 22627
rect 29779 22593 29788 22627
rect 29736 22584 29788 22593
rect 29828 22559 29880 22568
rect 29828 22525 29837 22559
rect 29837 22525 29871 22559
rect 29871 22525 29880 22559
rect 29828 22516 29880 22525
rect 29552 22448 29604 22500
rect 30380 22584 30432 22636
rect 31208 22584 31260 22636
rect 32864 22652 32916 22704
rect 32588 22627 32640 22636
rect 32588 22593 32597 22627
rect 32597 22593 32631 22627
rect 32631 22593 32640 22627
rect 32588 22584 32640 22593
rect 32772 22627 32824 22636
rect 32772 22593 32781 22627
rect 32781 22593 32815 22627
rect 32815 22593 32824 22627
rect 32772 22584 32824 22593
rect 36268 22627 36320 22636
rect 34244 22559 34296 22568
rect 34244 22525 34253 22559
rect 34253 22525 34287 22559
rect 34287 22525 34296 22559
rect 34244 22516 34296 22525
rect 34520 22516 34572 22568
rect 36268 22593 36277 22627
rect 36277 22593 36311 22627
rect 36311 22593 36320 22627
rect 36268 22584 36320 22593
rect 34612 22448 34664 22500
rect 16948 22380 17000 22432
rect 22284 22423 22336 22432
rect 22284 22389 22293 22423
rect 22293 22389 22327 22423
rect 22327 22389 22336 22423
rect 22284 22380 22336 22389
rect 22468 22380 22520 22432
rect 24216 22380 24268 22432
rect 30196 22423 30248 22432
rect 30196 22389 30205 22423
rect 30205 22389 30239 22423
rect 30239 22389 30248 22423
rect 30196 22380 30248 22389
rect 35624 22423 35676 22432
rect 35624 22389 35633 22423
rect 35633 22389 35667 22423
rect 35667 22389 35676 22423
rect 35624 22380 35676 22389
rect 37832 22423 37884 22432
rect 37832 22389 37841 22423
rect 37841 22389 37875 22423
rect 37875 22389 37884 22423
rect 37832 22380 37884 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 26792 22176 26844 22228
rect 28264 22219 28316 22228
rect 28264 22185 28273 22219
rect 28273 22185 28307 22219
rect 28307 22185 28316 22219
rect 28264 22176 28316 22185
rect 32588 22176 32640 22228
rect 34244 22176 34296 22228
rect 20720 22151 20772 22160
rect 20720 22117 20729 22151
rect 20729 22117 20763 22151
rect 20763 22117 20772 22151
rect 20720 22108 20772 22117
rect 1860 22083 1912 22092
rect 1860 22049 1869 22083
rect 1869 22049 1903 22083
rect 1903 22049 1912 22083
rect 1860 22040 1912 22049
rect 15752 22083 15804 22092
rect 15752 22049 15761 22083
rect 15761 22049 15795 22083
rect 15795 22049 15804 22083
rect 15752 22040 15804 22049
rect 16120 22040 16172 22092
rect 16488 22040 16540 22092
rect 20536 22040 20588 22092
rect 26700 22040 26752 22092
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 15660 22015 15712 22024
rect 15660 21981 15669 22015
rect 15669 21981 15703 22015
rect 15703 21981 15712 22015
rect 15660 21972 15712 21981
rect 15844 21972 15896 22024
rect 16580 22015 16632 22024
rect 16580 21981 16589 22015
rect 16589 21981 16623 22015
rect 16623 21981 16632 22015
rect 16580 21972 16632 21981
rect 16672 21972 16724 22024
rect 16948 22015 17000 22024
rect 16948 21981 16957 22015
rect 16957 21981 16991 22015
rect 16991 21981 17000 22015
rect 16948 21972 17000 21981
rect 20720 21972 20772 22024
rect 22376 22015 22428 22024
rect 22376 21981 22385 22015
rect 22385 21981 22419 22015
rect 22419 21981 22428 22015
rect 22376 21972 22428 21981
rect 22468 22015 22520 22024
rect 22468 21981 22477 22015
rect 22477 21981 22511 22015
rect 22511 21981 22520 22015
rect 22652 22015 22704 22024
rect 22468 21972 22520 21981
rect 22652 21981 22661 22015
rect 22661 21981 22695 22015
rect 22695 21981 22704 22015
rect 22652 21972 22704 21981
rect 23388 22015 23440 22024
rect 23388 21981 23397 22015
rect 23397 21981 23431 22015
rect 23431 21981 23440 22015
rect 23388 21972 23440 21981
rect 32128 22015 32180 22024
rect 2044 21904 2096 21956
rect 26424 21904 26476 21956
rect 32128 21981 32137 22015
rect 32137 21981 32171 22015
rect 32171 21981 32180 22015
rect 32128 21972 32180 21981
rect 32220 21972 32272 22024
rect 33692 21972 33744 22024
rect 34428 22040 34480 22092
rect 35532 22083 35584 22092
rect 35532 22049 35541 22083
rect 35541 22049 35575 22083
rect 35575 22049 35584 22083
rect 35532 22040 35584 22049
rect 37188 22083 37240 22092
rect 37188 22049 37197 22083
rect 37197 22049 37231 22083
rect 37231 22049 37240 22083
rect 37188 22040 37240 22049
rect 37832 22040 37884 22092
rect 34796 21972 34848 22024
rect 36268 21972 36320 22024
rect 37464 21904 37516 21956
rect 22560 21836 22612 21888
rect 27804 21836 27856 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 2044 21675 2096 21684
rect 2044 21641 2053 21675
rect 2053 21641 2087 21675
rect 2087 21641 2096 21675
rect 2044 21632 2096 21641
rect 16580 21632 16632 21684
rect 2412 21496 2464 21548
rect 15200 21564 15252 21616
rect 16212 21564 16264 21616
rect 18052 21632 18104 21684
rect 7840 21496 7892 21548
rect 8760 21471 8812 21480
rect 8760 21437 8769 21471
rect 8769 21437 8803 21471
rect 8803 21437 8812 21471
rect 8760 21428 8812 21437
rect 17500 21496 17552 21548
rect 19340 21564 19392 21616
rect 19616 21496 19668 21548
rect 19156 21428 19208 21480
rect 19984 21496 20036 21548
rect 20720 21632 20772 21684
rect 22652 21632 22704 21684
rect 26424 21675 26476 21684
rect 26424 21641 26433 21675
rect 26433 21641 26467 21675
rect 26467 21641 26476 21675
rect 26424 21632 26476 21641
rect 22284 21564 22336 21616
rect 22008 21539 22060 21548
rect 20352 21428 20404 21480
rect 22008 21505 22017 21539
rect 22017 21505 22051 21539
rect 22051 21505 22060 21539
rect 22008 21496 22060 21505
rect 22100 21496 22152 21548
rect 22560 21539 22612 21548
rect 22560 21505 22569 21539
rect 22569 21505 22603 21539
rect 22603 21505 22612 21539
rect 22560 21496 22612 21505
rect 24216 21539 24268 21548
rect 24216 21505 24234 21539
rect 24234 21505 24268 21539
rect 24216 21496 24268 21505
rect 25044 21539 25096 21548
rect 25044 21505 25053 21539
rect 25053 21505 25087 21539
rect 25087 21505 25096 21539
rect 25044 21496 25096 21505
rect 26424 21496 26476 21548
rect 26976 21539 27028 21548
rect 26976 21505 26985 21539
rect 26985 21505 27019 21539
rect 27019 21505 27028 21539
rect 26976 21496 27028 21505
rect 27804 21539 27856 21548
rect 17500 21360 17552 21412
rect 22468 21428 22520 21480
rect 26792 21428 26844 21480
rect 27804 21505 27813 21539
rect 27813 21505 27847 21539
rect 27847 21505 27856 21539
rect 27804 21496 27856 21505
rect 30472 21632 30524 21684
rect 32128 21675 32180 21684
rect 32128 21641 32137 21675
rect 32137 21641 32171 21675
rect 32171 21641 32180 21675
rect 32128 21632 32180 21641
rect 34520 21675 34572 21684
rect 34520 21641 34529 21675
rect 34529 21641 34563 21675
rect 34563 21641 34572 21675
rect 34520 21632 34572 21641
rect 30104 21496 30156 21548
rect 30380 21496 30432 21548
rect 31484 21496 31536 21548
rect 22928 21360 22980 21412
rect 26516 21292 26568 21344
rect 30840 21428 30892 21480
rect 33048 21496 33100 21548
rect 33324 21539 33376 21548
rect 33324 21505 33333 21539
rect 33333 21505 33367 21539
rect 33367 21505 33376 21539
rect 33324 21496 33376 21505
rect 34428 21539 34480 21548
rect 34428 21505 34437 21539
rect 34437 21505 34471 21539
rect 34471 21505 34480 21539
rect 34428 21496 34480 21505
rect 34796 21496 34848 21548
rect 35164 21496 35216 21548
rect 35624 21496 35676 21548
rect 36268 21632 36320 21684
rect 37464 21675 37516 21684
rect 37464 21641 37473 21675
rect 37473 21641 37507 21675
rect 37507 21641 37516 21675
rect 37464 21632 37516 21641
rect 30288 21360 30340 21412
rect 31208 21360 31260 21412
rect 32588 21428 32640 21480
rect 37648 21496 37700 21548
rect 37832 21428 37884 21480
rect 29092 21292 29144 21344
rect 31392 21292 31444 21344
rect 32772 21360 32824 21412
rect 33140 21292 33192 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1400 21088 1452 21140
rect 16120 21131 16172 21140
rect 16120 21097 16129 21131
rect 16129 21097 16163 21131
rect 16163 21097 16172 21131
rect 16120 21088 16172 21097
rect 16488 21088 16540 21140
rect 19984 21131 20036 21140
rect 19984 21097 19993 21131
rect 19993 21097 20027 21131
rect 20027 21097 20036 21131
rect 19984 21088 20036 21097
rect 26516 21131 26568 21140
rect 26516 21097 26525 21131
rect 26525 21097 26559 21131
rect 26559 21097 26568 21131
rect 26516 21088 26568 21097
rect 26976 21088 27028 21140
rect 29828 21088 29880 21140
rect 31944 21088 31996 21140
rect 8208 20995 8260 21004
rect 8208 20961 8217 20995
rect 8217 20961 8251 20995
rect 8251 20961 8260 20995
rect 8208 20952 8260 20961
rect 16212 20952 16264 21004
rect 7840 20884 7892 20936
rect 22652 20952 22704 21004
rect 23296 20995 23348 21004
rect 23296 20961 23305 20995
rect 23305 20961 23339 20995
rect 23339 20961 23348 20995
rect 23296 20952 23348 20961
rect 26700 20995 26752 21004
rect 26700 20961 26709 20995
rect 26709 20961 26743 20995
rect 26743 20961 26752 20995
rect 26700 20952 26752 20961
rect 30012 20952 30064 21004
rect 30380 20952 30432 21004
rect 31392 20995 31444 21004
rect 16672 20927 16724 20936
rect 16672 20893 16681 20927
rect 16681 20893 16715 20927
rect 16715 20893 16724 20927
rect 16672 20884 16724 20893
rect 20720 20884 20772 20936
rect 26424 20927 26476 20936
rect 26424 20893 26433 20927
rect 26433 20893 26467 20927
rect 26467 20893 26476 20927
rect 26424 20884 26476 20893
rect 17500 20816 17552 20868
rect 20352 20859 20404 20868
rect 20352 20825 20361 20859
rect 20361 20825 20395 20859
rect 20395 20825 20404 20859
rect 20352 20816 20404 20825
rect 26792 20816 26844 20868
rect 29920 20927 29972 20936
rect 29920 20893 29929 20927
rect 29929 20893 29963 20927
rect 29963 20893 29972 20927
rect 29920 20884 29972 20893
rect 29736 20816 29788 20868
rect 30288 20927 30340 20936
rect 30288 20893 30297 20927
rect 30297 20893 30331 20927
rect 30331 20893 30340 20927
rect 31392 20961 31401 20995
rect 31401 20961 31435 20995
rect 31435 20961 31444 20995
rect 31392 20952 31444 20961
rect 31484 20995 31536 21004
rect 31484 20961 31493 20995
rect 31493 20961 31527 20995
rect 31527 20961 31536 20995
rect 31484 20952 31536 20961
rect 30288 20884 30340 20893
rect 31208 20884 31260 20936
rect 26976 20748 27028 20800
rect 27160 20791 27212 20800
rect 27160 20757 27169 20791
rect 27169 20757 27203 20791
rect 27203 20757 27212 20791
rect 27160 20748 27212 20757
rect 30840 20748 30892 20800
rect 32588 20884 32640 20936
rect 32772 20927 32824 20936
rect 32772 20893 32781 20927
rect 32781 20893 32815 20927
rect 32815 20893 32824 20927
rect 34428 20952 34480 21004
rect 34520 20952 34572 21004
rect 33784 20927 33836 20936
rect 32772 20884 32824 20893
rect 33784 20893 33793 20927
rect 33793 20893 33827 20927
rect 33827 20893 33836 20927
rect 33784 20884 33836 20893
rect 33048 20816 33100 20868
rect 34060 20927 34112 20936
rect 34060 20893 34069 20927
rect 34069 20893 34103 20927
rect 34103 20893 34112 20927
rect 34060 20884 34112 20893
rect 34612 20884 34664 20936
rect 34796 20816 34848 20868
rect 31852 20748 31904 20800
rect 33692 20748 33744 20800
rect 38108 20995 38160 21004
rect 38108 20961 38117 20995
rect 38117 20961 38151 20995
rect 38151 20961 38160 20995
rect 38108 20952 38160 20961
rect 36268 20927 36320 20936
rect 36268 20893 36277 20927
rect 36277 20893 36311 20927
rect 36311 20893 36320 20927
rect 36268 20884 36320 20893
rect 35348 20791 35400 20800
rect 35348 20757 35357 20791
rect 35357 20757 35391 20791
rect 35391 20757 35400 20791
rect 35348 20748 35400 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 2320 20544 2372 20596
rect 7840 20476 7892 20528
rect 9220 20340 9272 20392
rect 26240 20544 26292 20596
rect 26424 20587 26476 20596
rect 26424 20553 26433 20587
rect 26433 20553 26467 20587
rect 26467 20553 26476 20587
rect 26424 20544 26476 20553
rect 29920 20544 29972 20596
rect 30012 20544 30064 20596
rect 33048 20587 33100 20596
rect 15752 20519 15804 20528
rect 15752 20485 15761 20519
rect 15761 20485 15795 20519
rect 15795 20485 15804 20519
rect 15752 20476 15804 20485
rect 16488 20476 16540 20528
rect 15660 20408 15712 20460
rect 15844 20451 15896 20460
rect 15844 20417 15853 20451
rect 15853 20417 15887 20451
rect 15887 20417 15896 20451
rect 22100 20476 22152 20528
rect 22836 20476 22888 20528
rect 15844 20408 15896 20417
rect 17500 20451 17552 20460
rect 17500 20417 17509 20451
rect 17509 20417 17543 20451
rect 17543 20417 17552 20451
rect 17500 20408 17552 20417
rect 18604 20340 18656 20392
rect 23296 20476 23348 20528
rect 30380 20476 30432 20528
rect 31668 20476 31720 20528
rect 33048 20553 33057 20587
rect 33057 20553 33091 20587
rect 33091 20553 33100 20587
rect 33048 20544 33100 20553
rect 33692 20587 33744 20596
rect 33692 20553 33701 20587
rect 33701 20553 33735 20587
rect 33735 20553 33744 20587
rect 33692 20544 33744 20553
rect 34060 20544 34112 20596
rect 23020 20408 23072 20460
rect 23388 20408 23440 20460
rect 25044 20451 25096 20460
rect 25044 20417 25053 20451
rect 25053 20417 25087 20451
rect 25087 20417 25096 20451
rect 25044 20408 25096 20417
rect 26976 20451 27028 20460
rect 26976 20417 26985 20451
rect 26985 20417 27019 20451
rect 27019 20417 27028 20451
rect 26976 20408 27028 20417
rect 27160 20451 27212 20460
rect 27160 20417 27169 20451
rect 27169 20417 27203 20451
rect 27203 20417 27212 20451
rect 27160 20408 27212 20417
rect 27896 20408 27948 20460
rect 29736 20408 29788 20460
rect 29920 20451 29972 20460
rect 29920 20417 29929 20451
rect 29929 20417 29963 20451
rect 29963 20417 29972 20451
rect 29920 20408 29972 20417
rect 29552 20340 29604 20392
rect 30196 20451 30248 20460
rect 30196 20417 30205 20451
rect 30205 20417 30239 20451
rect 30239 20417 30248 20451
rect 30932 20451 30984 20460
rect 30196 20408 30248 20417
rect 30932 20417 30941 20451
rect 30941 20417 30975 20451
rect 30975 20417 30984 20451
rect 30932 20408 30984 20417
rect 33140 20476 33192 20528
rect 34336 20408 34388 20460
rect 35532 20408 35584 20460
rect 36268 20408 36320 20460
rect 38200 20408 38252 20460
rect 23020 20272 23072 20324
rect 31760 20272 31812 20324
rect 33140 20340 33192 20392
rect 33692 20272 33744 20324
rect 34612 20315 34664 20324
rect 34612 20281 34621 20315
rect 34621 20281 34655 20315
rect 34655 20281 34664 20315
rect 34612 20272 34664 20281
rect 1400 20204 1452 20256
rect 15476 20204 15528 20256
rect 16856 20247 16908 20256
rect 16856 20213 16865 20247
rect 16865 20213 16899 20247
rect 16899 20213 16908 20247
rect 16856 20204 16908 20213
rect 17960 20204 18012 20256
rect 21824 20204 21876 20256
rect 22928 20247 22980 20256
rect 22928 20213 22937 20247
rect 22937 20213 22971 20247
rect 22971 20213 22980 20247
rect 22928 20204 22980 20213
rect 23572 20247 23624 20256
rect 23572 20213 23581 20247
rect 23581 20213 23615 20247
rect 23615 20213 23624 20247
rect 23572 20204 23624 20213
rect 26240 20204 26292 20256
rect 32496 20204 32548 20256
rect 37924 20204 37976 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 15752 20000 15804 20052
rect 15844 20000 15896 20052
rect 18052 20043 18104 20052
rect 18052 20009 18061 20043
rect 18061 20009 18095 20043
rect 18095 20009 18104 20043
rect 18052 20000 18104 20009
rect 20352 20000 20404 20052
rect 30288 20000 30340 20052
rect 30932 20000 30984 20052
rect 33324 20000 33376 20052
rect 23572 19932 23624 19984
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 1860 19907 1912 19916
rect 1860 19873 1869 19907
rect 1869 19873 1903 19907
rect 1903 19873 1912 19907
rect 1860 19864 1912 19873
rect 14188 19907 14240 19916
rect 14188 19873 14197 19907
rect 14197 19873 14231 19907
rect 14231 19873 14240 19907
rect 14188 19864 14240 19873
rect 18604 19864 18656 19916
rect 20168 19864 20220 19916
rect 22376 19864 22428 19916
rect 22836 19907 22888 19916
rect 22836 19873 22845 19907
rect 22845 19873 22879 19907
rect 22879 19873 22888 19907
rect 22836 19864 22888 19873
rect 26700 19864 26752 19916
rect 37188 19907 37240 19916
rect 37188 19873 37197 19907
rect 37197 19873 37231 19907
rect 37231 19873 37240 19907
rect 37188 19864 37240 19873
rect 37924 19907 37976 19916
rect 37924 19873 37933 19907
rect 37933 19873 37967 19907
rect 37967 19873 37976 19907
rect 37924 19864 37976 19873
rect 7840 19796 7892 19848
rect 17040 19796 17092 19848
rect 17868 19796 17920 19848
rect 20352 19839 20404 19848
rect 20352 19805 20361 19839
rect 20361 19805 20395 19839
rect 20395 19805 20404 19839
rect 20352 19796 20404 19805
rect 21824 19839 21876 19848
rect 1952 19728 2004 19780
rect 8116 19771 8168 19780
rect 8116 19737 8125 19771
rect 8125 19737 8159 19771
rect 8159 19737 8168 19771
rect 8116 19728 8168 19737
rect 15292 19728 15344 19780
rect 16856 19728 16908 19780
rect 17500 19728 17552 19780
rect 19432 19728 19484 19780
rect 19248 19660 19300 19712
rect 20076 19660 20128 19712
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 24952 19796 25004 19848
rect 26976 19796 27028 19848
rect 27620 19839 27672 19848
rect 27620 19805 27629 19839
rect 27629 19805 27663 19839
rect 27663 19805 27672 19839
rect 27620 19796 27672 19805
rect 24860 19771 24912 19780
rect 24860 19737 24869 19771
rect 24869 19737 24903 19771
rect 24903 19737 24912 19771
rect 24860 19728 24912 19737
rect 20904 19660 20956 19712
rect 24768 19660 24820 19712
rect 26148 19660 26200 19712
rect 28172 19796 28224 19848
rect 28908 19796 28960 19848
rect 30840 19839 30892 19848
rect 30840 19805 30849 19839
rect 30849 19805 30883 19839
rect 30883 19805 30892 19839
rect 30840 19796 30892 19805
rect 31668 19796 31720 19848
rect 33692 19796 33744 19848
rect 38108 19839 38160 19848
rect 38108 19805 38117 19839
rect 38117 19805 38151 19839
rect 38151 19805 38160 19839
rect 38108 19796 38160 19805
rect 27804 19660 27856 19712
rect 28264 19660 28316 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 2044 19363 2096 19372
rect 2044 19329 2053 19363
rect 2053 19329 2087 19363
rect 2087 19329 2096 19363
rect 16764 19456 16816 19508
rect 17960 19456 18012 19508
rect 19432 19456 19484 19508
rect 20352 19456 20404 19508
rect 22376 19456 22428 19508
rect 23388 19456 23440 19508
rect 26976 19499 27028 19508
rect 26976 19465 26985 19499
rect 26985 19465 27019 19499
rect 27019 19465 27028 19499
rect 26976 19456 27028 19465
rect 27620 19456 27672 19508
rect 28908 19456 28960 19508
rect 17868 19388 17920 19440
rect 15476 19363 15528 19372
rect 2044 19320 2096 19329
rect 15476 19329 15485 19363
rect 15485 19329 15519 19363
rect 15519 19329 15528 19363
rect 15476 19320 15528 19329
rect 15844 19320 15896 19372
rect 17960 19320 18012 19372
rect 19340 19320 19392 19372
rect 20996 19363 21048 19372
rect 22284 19388 22336 19440
rect 24768 19431 24820 19440
rect 24768 19397 24786 19431
rect 24786 19397 24820 19431
rect 24768 19388 24820 19397
rect 20996 19329 21014 19363
rect 21014 19329 21048 19363
rect 20996 19320 21048 19329
rect 22100 19363 22152 19372
rect 22100 19329 22134 19363
rect 22134 19329 22152 19363
rect 25044 19363 25096 19372
rect 22100 19320 22152 19329
rect 25044 19329 25053 19363
rect 25053 19329 25087 19363
rect 25087 19329 25096 19363
rect 25044 19320 25096 19329
rect 26148 19320 26200 19372
rect 27160 19363 27212 19372
rect 27160 19329 27169 19363
rect 27169 19329 27203 19363
rect 27203 19329 27212 19363
rect 27160 19320 27212 19329
rect 28540 19388 28592 19440
rect 28264 19363 28316 19372
rect 28264 19329 28298 19363
rect 28298 19329 28316 19363
rect 28264 19320 28316 19329
rect 33140 19320 33192 19372
rect 34244 19320 34296 19372
rect 38108 19320 38160 19372
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 15752 19295 15804 19304
rect 15752 19261 15761 19295
rect 15761 19261 15795 19295
rect 15795 19261 15804 19295
rect 15752 19252 15804 19261
rect 18144 19252 18196 19304
rect 27896 19252 27948 19304
rect 33784 19252 33836 19304
rect 34336 19295 34388 19304
rect 34336 19261 34345 19295
rect 34345 19261 34379 19295
rect 34379 19261 34388 19295
rect 34336 19252 34388 19261
rect 26608 19116 26660 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 17960 18912 18012 18964
rect 19248 18912 19300 18964
rect 19340 18912 19392 18964
rect 20996 18912 21048 18964
rect 22100 18955 22152 18964
rect 22100 18921 22109 18955
rect 22109 18921 22143 18955
rect 22143 18921 22152 18955
rect 22100 18912 22152 18921
rect 22836 18912 22888 18964
rect 24860 18912 24912 18964
rect 27896 18955 27948 18964
rect 27896 18921 27905 18955
rect 27905 18921 27939 18955
rect 27939 18921 27948 18955
rect 27896 18912 27948 18921
rect 28172 18912 28224 18964
rect 18144 18776 18196 18828
rect 18052 18708 18104 18760
rect 20352 18776 20404 18828
rect 19248 18751 19300 18760
rect 19248 18717 19257 18751
rect 19257 18717 19291 18751
rect 19291 18717 19300 18751
rect 19248 18708 19300 18717
rect 19340 18708 19392 18760
rect 20076 18751 20128 18760
rect 20076 18717 20085 18751
rect 20085 18717 20119 18751
rect 20119 18717 20128 18751
rect 20076 18708 20128 18717
rect 20904 18751 20956 18760
rect 19984 18640 20036 18692
rect 20904 18717 20913 18751
rect 20913 18717 20947 18751
rect 20947 18717 20956 18751
rect 20904 18708 20956 18717
rect 27252 18776 27304 18828
rect 17316 18572 17368 18624
rect 22836 18708 22888 18760
rect 26608 18751 26660 18760
rect 26608 18717 26617 18751
rect 26617 18717 26651 18751
rect 26651 18717 26660 18751
rect 26608 18708 26660 18717
rect 26792 18751 26844 18760
rect 26792 18717 26801 18751
rect 26801 18717 26835 18751
rect 26835 18717 26844 18751
rect 26792 18708 26844 18717
rect 31760 18819 31812 18828
rect 31760 18785 31769 18819
rect 31769 18785 31803 18819
rect 31803 18785 31812 18819
rect 31760 18776 31812 18785
rect 23020 18683 23072 18692
rect 23020 18649 23029 18683
rect 23029 18649 23063 18683
rect 23063 18649 23072 18683
rect 23020 18640 23072 18649
rect 27620 18640 27672 18692
rect 29092 18640 29144 18692
rect 30840 18751 30892 18760
rect 30840 18717 30849 18751
rect 30849 18717 30883 18751
rect 30883 18717 30892 18751
rect 30840 18708 30892 18717
rect 31852 18751 31904 18760
rect 30104 18640 30156 18692
rect 31852 18717 31861 18751
rect 31861 18717 31895 18751
rect 31895 18717 31904 18751
rect 31852 18708 31904 18717
rect 33140 18776 33192 18828
rect 35348 18776 35400 18828
rect 32312 18640 32364 18692
rect 33784 18708 33836 18760
rect 36268 18751 36320 18760
rect 36268 18717 36277 18751
rect 36277 18717 36311 18751
rect 36311 18717 36320 18751
rect 36268 18708 36320 18717
rect 36452 18683 36504 18692
rect 36452 18649 36461 18683
rect 36461 18649 36495 18683
rect 36495 18649 36504 18683
rect 36452 18640 36504 18649
rect 38108 18683 38160 18692
rect 38108 18649 38117 18683
rect 38117 18649 38151 18683
rect 38151 18649 38160 18683
rect 38108 18640 38160 18649
rect 23296 18572 23348 18624
rect 26424 18615 26476 18624
rect 26424 18581 26433 18615
rect 26433 18581 26467 18615
rect 26467 18581 26476 18615
rect 26424 18572 26476 18581
rect 26792 18572 26844 18624
rect 27160 18572 27212 18624
rect 28540 18615 28592 18624
rect 28540 18581 28549 18615
rect 28549 18581 28583 18615
rect 28583 18581 28592 18615
rect 28540 18572 28592 18581
rect 31300 18572 31352 18624
rect 31576 18572 31628 18624
rect 32956 18615 33008 18624
rect 32956 18581 32965 18615
rect 32965 18581 32999 18615
rect 32999 18581 33008 18615
rect 32956 18572 33008 18581
rect 34704 18615 34756 18624
rect 34704 18581 34713 18615
rect 34713 18581 34747 18615
rect 34747 18581 34756 18615
rect 34704 18572 34756 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 18144 18368 18196 18420
rect 19340 18411 19392 18420
rect 19340 18377 19349 18411
rect 19349 18377 19383 18411
rect 19383 18377 19392 18411
rect 19340 18368 19392 18377
rect 30104 18368 30156 18420
rect 32220 18368 32272 18420
rect 33140 18368 33192 18420
rect 34244 18368 34296 18420
rect 36452 18368 36504 18420
rect 7380 18300 7432 18352
rect 8116 18300 8168 18352
rect 17040 18275 17092 18284
rect 17040 18241 17049 18275
rect 17049 18241 17083 18275
rect 17083 18241 17092 18275
rect 17040 18232 17092 18241
rect 17316 18275 17368 18284
rect 17316 18241 17350 18275
rect 17350 18241 17368 18275
rect 17316 18232 17368 18241
rect 19432 18232 19484 18284
rect 28448 18275 28500 18284
rect 28448 18241 28457 18275
rect 28457 18241 28491 18275
rect 28491 18241 28500 18275
rect 28448 18232 28500 18241
rect 28540 18232 28592 18284
rect 31300 18275 31352 18284
rect 31300 18241 31309 18275
rect 31309 18241 31343 18275
rect 31343 18241 31352 18275
rect 31300 18232 31352 18241
rect 31576 18275 31628 18284
rect 31576 18241 31585 18275
rect 31585 18241 31619 18275
rect 31619 18241 31628 18275
rect 31576 18232 31628 18241
rect 32680 18232 32732 18284
rect 33232 18275 33284 18284
rect 33232 18241 33266 18275
rect 33266 18241 33284 18275
rect 33232 18232 33284 18241
rect 36268 18232 36320 18284
rect 37464 18275 37516 18284
rect 37464 18241 37473 18275
rect 37473 18241 37507 18275
rect 37507 18241 37516 18275
rect 37464 18232 37516 18241
rect 19984 18164 20036 18216
rect 31116 18164 31168 18216
rect 32772 18164 32824 18216
rect 20168 18096 20220 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 31208 18071 31260 18080
rect 31208 18037 31217 18071
rect 31217 18037 31251 18071
rect 31251 18037 31260 18071
rect 31208 18028 31260 18037
rect 36084 18071 36136 18080
rect 36084 18037 36093 18071
rect 36093 18037 36127 18071
rect 36127 18037 36136 18071
rect 36084 18028 36136 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 27252 17824 27304 17876
rect 30840 17824 30892 17876
rect 32956 17824 33008 17876
rect 33232 17756 33284 17808
rect 1676 17688 1728 17740
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 25044 17688 25096 17740
rect 32680 17688 32732 17740
rect 32772 17688 32824 17740
rect 36084 17688 36136 17740
rect 38108 17731 38160 17740
rect 38108 17697 38117 17731
rect 38117 17697 38151 17731
rect 38151 17697 38160 17731
rect 38108 17688 38160 17697
rect 26424 17620 26476 17672
rect 33140 17663 33192 17672
rect 33140 17629 33149 17663
rect 33149 17629 33183 17663
rect 33183 17629 33192 17663
rect 33140 17620 33192 17629
rect 34704 17620 34756 17672
rect 2136 17552 2188 17604
rect 31208 17552 31260 17604
rect 36452 17595 36504 17604
rect 36452 17561 36461 17595
rect 36461 17561 36495 17595
rect 36495 17561 36504 17595
rect 36452 17552 36504 17561
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 2136 17323 2188 17332
rect 2136 17289 2145 17323
rect 2145 17289 2179 17323
rect 2179 17289 2188 17323
rect 2136 17280 2188 17289
rect 36452 17280 36504 17332
rect 2228 17187 2280 17196
rect 2228 17153 2237 17187
rect 2237 17153 2271 17187
rect 2271 17153 2280 17187
rect 2228 17144 2280 17153
rect 15384 17144 15436 17196
rect 15568 17144 15620 17196
rect 37464 17187 37516 17196
rect 37464 17153 37473 17187
rect 37473 17153 37507 17187
rect 37507 17153 37516 17187
rect 37464 17144 37516 17153
rect 37648 17144 37700 17196
rect 1400 16983 1452 16992
rect 1400 16949 1409 16983
rect 1409 16949 1443 16983
rect 1443 16949 1452 16983
rect 1400 16940 1452 16949
rect 36268 16940 36320 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1400 16643 1452 16652
rect 1400 16609 1409 16643
rect 1409 16609 1443 16643
rect 1443 16609 1452 16643
rect 1400 16600 1452 16609
rect 1860 16643 1912 16652
rect 1860 16609 1869 16643
rect 1869 16609 1903 16643
rect 1903 16609 1912 16643
rect 1860 16600 1912 16609
rect 36268 16643 36320 16652
rect 36268 16609 36277 16643
rect 36277 16609 36311 16643
rect 36311 16609 36320 16643
rect 36268 16600 36320 16609
rect 38108 16643 38160 16652
rect 38108 16609 38117 16643
rect 38117 16609 38151 16643
rect 38151 16609 38160 16643
rect 38108 16600 38160 16609
rect 2044 16464 2096 16516
rect 36452 16507 36504 16516
rect 36452 16473 36461 16507
rect 36461 16473 36495 16507
rect 36495 16473 36504 16507
rect 36452 16464 36504 16473
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2044 16235 2096 16244
rect 2044 16201 2053 16235
rect 2053 16201 2087 16235
rect 2087 16201 2096 16235
rect 2044 16192 2096 16201
rect 36452 16192 36504 16244
rect 2136 16099 2188 16108
rect 2136 16065 2145 16099
rect 2145 16065 2179 16099
rect 2179 16065 2188 16099
rect 2136 16056 2188 16065
rect 37464 16099 37516 16108
rect 37464 16065 37473 16099
rect 37473 16065 37507 16099
rect 37507 16065 37516 16099
rect 37464 16056 37516 16065
rect 38016 16056 38068 16108
rect 3240 15852 3292 15904
rect 36268 15852 36320 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1400 15555 1452 15564
rect 1400 15521 1409 15555
rect 1409 15521 1443 15555
rect 1443 15521 1452 15555
rect 1400 15512 1452 15521
rect 3240 15555 3292 15564
rect 3240 15521 3249 15555
rect 3249 15521 3283 15555
rect 3283 15521 3292 15555
rect 3240 15512 3292 15521
rect 36268 15555 36320 15564
rect 36268 15521 36277 15555
rect 36277 15521 36311 15555
rect 36311 15521 36320 15555
rect 36268 15512 36320 15521
rect 38108 15555 38160 15564
rect 38108 15521 38117 15555
rect 38117 15521 38151 15555
rect 38151 15521 38160 15555
rect 38108 15512 38160 15521
rect 3056 15419 3108 15428
rect 3056 15385 3065 15419
rect 3065 15385 3099 15419
rect 3099 15385 3108 15419
rect 3056 15376 3108 15385
rect 36452 15419 36504 15428
rect 36452 15385 36461 15419
rect 36461 15385 36495 15419
rect 36495 15385 36504 15419
rect 36452 15376 36504 15385
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 3056 15104 3108 15156
rect 36452 15104 36504 15156
rect 2320 14968 2372 15020
rect 14464 14968 14516 15020
rect 36360 14968 36412 15020
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1676 14356 1728 14408
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1860 13472 1912 13524
rect 1676 13268 1728 13320
rect 2228 13311 2280 13320
rect 2228 13277 2237 13311
rect 2237 13277 2271 13311
rect 2271 13277 2280 13311
rect 2228 13268 2280 13277
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 37832 12903 37884 12912
rect 37832 12869 37841 12903
rect 37841 12869 37875 12903
rect 37875 12869 37884 12903
rect 37832 12860 37884 12869
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 38108 12835 38160 12844
rect 38108 12801 38117 12835
rect 38117 12801 38151 12835
rect 38151 12801 38160 12835
rect 38108 12792 38160 12801
rect 1860 12767 1912 12776
rect 1860 12733 1869 12767
rect 1869 12733 1903 12767
rect 1903 12733 1912 12767
rect 1860 12724 1912 12733
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1860 12384 1912 12436
rect 9404 12180 9456 12232
rect 38108 12180 38160 12232
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 8760 11704 8812 11756
rect 37372 11747 37424 11756
rect 37372 11713 37381 11747
rect 37381 11713 37415 11747
rect 37415 11713 37424 11747
rect 37372 11704 37424 11713
rect 37924 11500 37976 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 37188 11203 37240 11212
rect 37188 11169 37197 11203
rect 37197 11169 37231 11203
rect 37231 11169 37240 11203
rect 37188 11160 37240 11169
rect 37924 11203 37976 11212
rect 37924 11169 37933 11203
rect 37933 11169 37967 11203
rect 37967 11169 37976 11203
rect 37924 11160 37976 11169
rect 38108 11203 38160 11212
rect 38108 11169 38117 11203
rect 38117 11169 38151 11203
rect 38151 11169 38160 11203
rect 38108 11160 38160 11169
rect 2136 11092 2188 11144
rect 3424 11092 3476 11144
rect 3240 11024 3292 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 3240 10727 3292 10736
rect 3240 10693 3249 10727
rect 3249 10693 3283 10727
rect 3283 10693 3292 10727
rect 3240 10684 3292 10693
rect 3424 10659 3476 10668
rect 3424 10625 3433 10659
rect 3433 10625 3467 10659
rect 3467 10625 3476 10659
rect 3424 10616 3476 10625
rect 37556 10616 37608 10668
rect 1584 10591 1636 10600
rect 1584 10557 1593 10591
rect 1593 10557 1627 10591
rect 1627 10557 1636 10591
rect 1584 10548 1636 10557
rect 36452 10412 36504 10464
rect 38108 10455 38160 10464
rect 38108 10421 38117 10455
rect 38117 10421 38151 10455
rect 38151 10421 38160 10455
rect 38108 10412 38160 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 36452 10115 36504 10124
rect 36452 10081 36461 10115
rect 36461 10081 36495 10115
rect 36495 10081 36504 10115
rect 36452 10072 36504 10081
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 20352 10004 20404 10056
rect 36268 10047 36320 10056
rect 36268 10013 36277 10047
rect 36277 10013 36311 10047
rect 36311 10013 36320 10047
rect 36268 10004 36320 10013
rect 38016 9936 38068 9988
rect 2044 9868 2096 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2044 9639 2096 9648
rect 2044 9605 2053 9639
rect 2053 9605 2087 9639
rect 2087 9605 2096 9639
rect 2044 9596 2096 9605
rect 1860 9571 1912 9580
rect 1860 9537 1869 9571
rect 1869 9537 1903 9571
rect 1903 9537 1912 9571
rect 1860 9528 1912 9537
rect 36268 9528 36320 9580
rect 37464 9571 37516 9580
rect 37464 9537 37473 9571
rect 37473 9537 37507 9571
rect 37507 9537 37516 9571
rect 37464 9528 37516 9537
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 37924 9324 37976 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 37188 9027 37240 9036
rect 37188 8993 37197 9027
rect 37197 8993 37231 9027
rect 37231 8993 37240 9027
rect 37188 8984 37240 8993
rect 37924 9027 37976 9036
rect 37924 8993 37933 9027
rect 37933 8993 37967 9027
rect 37967 8993 37976 9027
rect 37924 8984 37976 8993
rect 38108 9027 38160 9036
rect 38108 8993 38117 9027
rect 38117 8993 38151 9027
rect 38151 8993 38160 9027
rect 38108 8984 38160 8993
rect 2044 8959 2096 8968
rect 2044 8925 2053 8959
rect 2053 8925 2087 8959
rect 2087 8925 2096 8959
rect 2044 8916 2096 8925
rect 2872 8916 2924 8968
rect 2228 8780 2280 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 2228 8551 2280 8560
rect 2228 8517 2237 8551
rect 2237 8517 2271 8551
rect 2271 8517 2280 8551
rect 2228 8508 2280 8517
rect 2044 8483 2096 8492
rect 2044 8449 2053 8483
rect 2053 8449 2087 8483
rect 2087 8449 2096 8483
rect 2044 8440 2096 8449
rect 2872 8415 2924 8424
rect 2872 8381 2881 8415
rect 2881 8381 2915 8415
rect 2915 8381 2924 8415
rect 2872 8372 2924 8381
rect 38108 8304 38160 8356
rect 1400 8279 1452 8288
rect 1400 8245 1409 8279
rect 1409 8245 1443 8279
rect 1443 8245 1452 8279
rect 1400 8236 1452 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 1400 7939 1452 7948
rect 1400 7905 1409 7939
rect 1409 7905 1443 7939
rect 1443 7905 1452 7939
rect 1400 7896 1452 7905
rect 2780 7939 2832 7948
rect 2780 7905 2789 7939
rect 2789 7905 2823 7939
rect 2823 7905 2832 7939
rect 2780 7896 2832 7905
rect 37832 7871 37884 7880
rect 37832 7837 37841 7871
rect 37841 7837 37875 7871
rect 37875 7837 37884 7871
rect 37832 7828 37884 7837
rect 2228 7760 2280 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2228 7531 2280 7540
rect 2228 7497 2237 7531
rect 2237 7497 2271 7531
rect 2271 7497 2280 7531
rect 2228 7488 2280 7497
rect 7012 7352 7064 7404
rect 37648 7352 37700 7404
rect 1400 7148 1452 7200
rect 37924 7148 37976 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1400 6851 1452 6860
rect 1400 6817 1409 6851
rect 1409 6817 1443 6851
rect 1443 6817 1452 6851
rect 1400 6808 1452 6817
rect 2780 6851 2832 6860
rect 2780 6817 2789 6851
rect 2789 6817 2823 6851
rect 2823 6817 2832 6851
rect 37188 6851 37240 6860
rect 2780 6808 2832 6817
rect 37188 6817 37197 6851
rect 37197 6817 37231 6851
rect 37231 6817 37240 6851
rect 37188 6808 37240 6817
rect 37924 6851 37976 6860
rect 37924 6817 37933 6851
rect 37933 6817 37967 6851
rect 37967 6817 37976 6851
rect 37924 6808 37976 6817
rect 38108 6851 38160 6860
rect 38108 6817 38117 6851
rect 38117 6817 38151 6851
rect 38151 6817 38160 6851
rect 38108 6808 38160 6817
rect 2044 6672 2096 6724
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2044 6443 2096 6452
rect 2044 6409 2053 6443
rect 2053 6409 2087 6443
rect 2087 6409 2096 6443
rect 2044 6400 2096 6409
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 2412 6264 2464 6316
rect 37556 6264 37608 6316
rect 35348 6239 35400 6248
rect 35348 6205 35357 6239
rect 35357 6205 35391 6239
rect 35391 6205 35400 6239
rect 35348 6196 35400 6205
rect 36544 6239 36596 6248
rect 36544 6205 36553 6239
rect 36553 6205 36587 6239
rect 36587 6205 36596 6239
rect 36544 6196 36596 6205
rect 37832 6196 37884 6248
rect 3240 6060 3292 6112
rect 37924 6060 37976 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 37740 5788 37792 5840
rect 3240 5763 3292 5772
rect 3240 5729 3249 5763
rect 3249 5729 3283 5763
rect 3283 5729 3292 5763
rect 3240 5720 3292 5729
rect 37188 5763 37240 5772
rect 37188 5729 37197 5763
rect 37197 5729 37231 5763
rect 37231 5729 37240 5763
rect 37188 5720 37240 5729
rect 37924 5763 37976 5772
rect 37924 5729 37933 5763
rect 37933 5729 37967 5763
rect 37967 5729 37976 5763
rect 37924 5720 37976 5729
rect 33416 5695 33468 5704
rect 33416 5661 33425 5695
rect 33425 5661 33459 5695
rect 33459 5661 33468 5695
rect 33416 5652 33468 5661
rect 34520 5652 34572 5704
rect 36452 5652 36504 5704
rect 1400 5627 1452 5636
rect 1400 5593 1409 5627
rect 1409 5593 1443 5627
rect 1443 5593 1452 5627
rect 1400 5584 1452 5593
rect 3056 5627 3108 5636
rect 3056 5593 3065 5627
rect 3065 5593 3099 5627
rect 3099 5593 3108 5627
rect 3056 5584 3108 5593
rect 35532 5516 35584 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3056 5312 3108 5364
rect 36544 5312 36596 5364
rect 14556 5244 14608 5296
rect 35256 5287 35308 5296
rect 2320 5176 2372 5228
rect 32680 5219 32732 5228
rect 32680 5185 32689 5219
rect 32689 5185 32723 5219
rect 32723 5185 32732 5219
rect 32680 5176 32732 5185
rect 33416 5219 33468 5228
rect 33416 5185 33425 5219
rect 33425 5185 33459 5219
rect 33459 5185 33468 5219
rect 33416 5176 33468 5185
rect 35256 5253 35265 5287
rect 35265 5253 35299 5287
rect 35299 5253 35308 5287
rect 35256 5244 35308 5253
rect 37832 5176 37884 5228
rect 2964 5151 3016 5160
rect 2964 5117 2973 5151
rect 2973 5117 3007 5151
rect 3007 5117 3016 5151
rect 2964 5108 3016 5117
rect 3884 5108 3936 5160
rect 3976 5151 4028 5160
rect 3976 5117 3985 5151
rect 3985 5117 4019 5151
rect 4019 5117 4028 5151
rect 3976 5108 4028 5117
rect 33968 5040 34020 5092
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 8944 4972 8996 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2964 4811 3016 4820
rect 2964 4777 2973 4811
rect 2973 4777 3007 4811
rect 3007 4777 3016 4811
rect 2964 4768 3016 4777
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 4068 4700 4120 4752
rect 6184 4632 6236 4684
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 15476 4632 15528 4684
rect 34612 4700 34664 4752
rect 33968 4675 34020 4684
rect 33968 4641 33977 4675
rect 33977 4641 34011 4675
rect 34011 4641 34020 4675
rect 33968 4632 34020 4641
rect 34520 4632 34572 4684
rect 35532 4675 35584 4684
rect 35532 4641 35541 4675
rect 35541 4641 35575 4675
rect 35575 4641 35584 4675
rect 35532 4632 35584 4641
rect 36084 4675 36136 4684
rect 36084 4641 36093 4675
rect 36093 4641 36127 4675
rect 36127 4641 36136 4675
rect 36084 4632 36136 4641
rect 1400 4564 1452 4616
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 8208 4564 8260 4616
rect 9864 4607 9916 4616
rect 9864 4573 9873 4607
rect 9873 4573 9907 4607
rect 9907 4573 9916 4607
rect 9864 4564 9916 4573
rect 15200 4607 15252 4616
rect 15200 4573 15209 4607
rect 15209 4573 15243 4607
rect 15243 4573 15252 4607
rect 15200 4564 15252 4573
rect 24400 4564 24452 4616
rect 37372 4564 37424 4616
rect 5816 4496 5868 4548
rect 7288 4496 7340 4548
rect 15384 4539 15436 4548
rect 15384 4505 15393 4539
rect 15393 4505 15427 4539
rect 15427 4505 15436 4539
rect 15384 4496 15436 4505
rect 9312 4471 9364 4480
rect 9312 4437 9321 4471
rect 9321 4437 9355 4471
rect 9355 4437 9364 4471
rect 9312 4428 9364 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 3976 4224 4028 4276
rect 9496 4156 9548 4208
rect 15384 4224 15436 4276
rect 4712 4131 4764 4140
rect 4712 4097 4721 4131
rect 4721 4097 4755 4131
rect 4755 4097 4764 4131
rect 4712 4088 4764 4097
rect 7104 4088 7156 4140
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 1952 4063 2004 4072
rect 1952 4029 1961 4063
rect 1961 4029 1995 4063
rect 1995 4029 2004 4063
rect 1952 4020 2004 4029
rect 2504 4020 2556 4072
rect 8668 4063 8720 4072
rect 664 3952 716 4004
rect 8668 4029 8677 4063
rect 8677 4029 8711 4063
rect 8711 4029 8720 4063
rect 8668 4020 8720 4029
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 6552 3884 6604 3936
rect 6644 3884 6696 3936
rect 9404 4020 9456 4072
rect 9496 3952 9548 4004
rect 15752 4156 15804 4208
rect 23664 4156 23716 4208
rect 15660 4131 15712 4140
rect 15660 4097 15669 4131
rect 15669 4097 15703 4131
rect 15703 4097 15712 4131
rect 15660 4088 15712 4097
rect 20352 4131 20404 4140
rect 20352 4097 20361 4131
rect 20361 4097 20395 4131
rect 20395 4097 20404 4131
rect 20352 4088 20404 4097
rect 22192 4131 22244 4140
rect 22192 4097 22201 4131
rect 22201 4097 22235 4131
rect 22235 4097 22244 4131
rect 22192 4088 22244 4097
rect 32220 4131 32272 4140
rect 32220 4097 32229 4131
rect 32229 4097 32263 4131
rect 32263 4097 32272 4131
rect 32220 4088 32272 4097
rect 37280 4088 37332 4140
rect 22560 4020 22612 4072
rect 23572 4063 23624 4072
rect 23572 4029 23581 4063
rect 23581 4029 23615 4063
rect 23615 4029 23624 4063
rect 23572 4020 23624 4029
rect 23848 4063 23900 4072
rect 23848 4029 23857 4063
rect 23857 4029 23891 4063
rect 23891 4029 23900 4063
rect 23848 4020 23900 4029
rect 32496 4063 32548 4072
rect 32496 4029 32505 4063
rect 32505 4029 32539 4063
rect 32539 4029 32548 4063
rect 32496 4020 32548 4029
rect 34152 4020 34204 4072
rect 34980 4063 35032 4072
rect 34980 4029 34989 4063
rect 34989 4029 35023 4063
rect 35023 4029 35032 4063
rect 34980 4020 35032 4029
rect 35440 4063 35492 4072
rect 35440 4029 35449 4063
rect 35449 4029 35483 4063
rect 35483 4029 35492 4063
rect 35440 4020 35492 4029
rect 13820 3952 13872 4004
rect 14832 3952 14884 4004
rect 10416 3884 10468 3936
rect 11888 3884 11940 3936
rect 18144 3927 18196 3936
rect 18144 3893 18153 3927
rect 18153 3893 18187 3927
rect 18187 3893 18196 3927
rect 18144 3884 18196 3893
rect 20168 3884 20220 3936
rect 24584 3884 24636 3936
rect 37280 3884 37332 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2504 3723 2556 3732
rect 2504 3689 2513 3723
rect 2513 3689 2547 3723
rect 2547 3689 2556 3723
rect 2504 3680 2556 3689
rect 2136 3476 2188 3528
rect 5356 3612 5408 3664
rect 8668 3680 8720 3732
rect 32496 3680 32548 3732
rect 34152 3723 34204 3732
rect 34152 3689 34161 3723
rect 34161 3689 34195 3723
rect 34195 3689 34204 3723
rect 34152 3680 34204 3689
rect 34796 3680 34848 3732
rect 15200 3612 15252 3664
rect 22560 3655 22612 3664
rect 4804 3587 4856 3596
rect 4804 3553 4813 3587
rect 4813 3553 4847 3587
rect 4847 3553 4856 3587
rect 4804 3544 4856 3553
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 2964 3408 3016 3460
rect 7012 3476 7064 3528
rect 10232 3544 10284 3596
rect 10416 3587 10468 3596
rect 10416 3553 10425 3587
rect 10425 3553 10459 3587
rect 10459 3553 10468 3587
rect 10416 3544 10468 3553
rect 10968 3587 11020 3596
rect 10968 3553 10977 3587
rect 10977 3553 11011 3587
rect 11011 3553 11020 3587
rect 10968 3544 11020 3553
rect 16764 3587 16816 3596
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 1584 3340 1636 3392
rect 3148 3383 3200 3392
rect 3148 3349 3157 3383
rect 3157 3349 3191 3383
rect 3191 3349 3200 3383
rect 3148 3340 3200 3349
rect 6828 3340 6880 3392
rect 9128 3340 9180 3392
rect 16764 3553 16773 3587
rect 16773 3553 16807 3587
rect 16807 3553 16816 3587
rect 16764 3544 16816 3553
rect 15568 3519 15620 3528
rect 11704 3340 11756 3392
rect 15568 3485 15577 3519
rect 15577 3485 15611 3519
rect 15611 3485 15620 3519
rect 15568 3476 15620 3485
rect 16212 3519 16264 3528
rect 16212 3485 16221 3519
rect 16221 3485 16255 3519
rect 16255 3485 16264 3519
rect 16212 3476 16264 3485
rect 22560 3621 22569 3655
rect 22569 3621 22603 3655
rect 22603 3621 22612 3655
rect 22560 3612 22612 3621
rect 23572 3612 23624 3664
rect 20168 3587 20220 3596
rect 20168 3553 20177 3587
rect 20177 3553 20211 3587
rect 20211 3553 20220 3587
rect 20168 3544 20220 3553
rect 20628 3587 20680 3596
rect 20628 3553 20637 3587
rect 20637 3553 20671 3587
rect 20671 3553 20680 3587
rect 20628 3544 20680 3553
rect 24400 3587 24452 3596
rect 24400 3553 24409 3587
rect 24409 3553 24443 3587
rect 24443 3553 24452 3587
rect 24400 3544 24452 3553
rect 24584 3587 24636 3596
rect 24584 3553 24593 3587
rect 24593 3553 24627 3587
rect 24627 3553 24636 3587
rect 24584 3544 24636 3553
rect 18788 3476 18840 3528
rect 22560 3476 22612 3528
rect 23020 3519 23072 3528
rect 23020 3485 23029 3519
rect 23029 3485 23063 3519
rect 23063 3485 23072 3519
rect 23020 3476 23072 3485
rect 23664 3519 23716 3528
rect 23664 3485 23673 3519
rect 23673 3485 23707 3519
rect 23707 3485 23716 3519
rect 23664 3476 23716 3485
rect 24124 3476 24176 3528
rect 32220 3544 32272 3596
rect 18328 3340 18380 3392
rect 24032 3340 24084 3392
rect 24124 3340 24176 3392
rect 27804 3408 27856 3460
rect 32588 3476 32640 3528
rect 33232 3476 33284 3528
rect 37464 3544 37516 3596
rect 35624 3519 35676 3528
rect 35624 3485 35633 3519
rect 35633 3485 35667 3519
rect 35667 3485 35676 3519
rect 35624 3476 35676 3485
rect 38108 3519 38160 3528
rect 38108 3485 38117 3519
rect 38117 3485 38151 3519
rect 38151 3485 38160 3519
rect 38108 3476 38160 3485
rect 35808 3408 35860 3460
rect 37464 3408 37516 3460
rect 27988 3340 28040 3392
rect 33416 3340 33468 3392
rect 35716 3383 35768 3392
rect 35716 3349 35725 3383
rect 35725 3349 35759 3383
rect 35759 3349 35768 3383
rect 35716 3340 35768 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 3148 3111 3200 3120
rect 3148 3077 3157 3111
rect 3157 3077 3191 3111
rect 3191 3077 3200 3111
rect 3148 3068 3200 3077
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2964 3043 3016 3052
rect 2964 3009 2973 3043
rect 2973 3009 3007 3043
rect 3007 3009 3016 3043
rect 2964 3000 3016 3009
rect 6828 3111 6880 3120
rect 6828 3077 6837 3111
rect 6837 3077 6871 3111
rect 6871 3077 6880 3111
rect 6828 3068 6880 3077
rect 7104 3136 7156 3188
rect 13820 3136 13872 3188
rect 15660 3136 15712 3188
rect 8300 3068 8352 3120
rect 9128 3111 9180 3120
rect 9128 3077 9137 3111
rect 9137 3077 9171 3111
rect 9171 3077 9180 3111
rect 9128 3068 9180 3077
rect 11888 3111 11940 3120
rect 11888 3077 11897 3111
rect 11897 3077 11931 3111
rect 11931 3077 11940 3111
rect 11888 3068 11940 3077
rect 18328 3111 18380 3120
rect 18328 3077 18337 3111
rect 18337 3077 18371 3111
rect 18371 3077 18380 3111
rect 18328 3068 18380 3077
rect 24032 3111 24084 3120
rect 24032 3077 24041 3111
rect 24041 3077 24075 3111
rect 24075 3077 24084 3111
rect 24032 3068 24084 3077
rect 27988 3111 28040 3120
rect 27988 3077 27997 3111
rect 27997 3077 28031 3111
rect 28031 3077 28040 3111
rect 27988 3068 28040 3077
rect 33416 3111 33468 3120
rect 33416 3077 33425 3111
rect 33425 3077 33459 3111
rect 33459 3077 33468 3111
rect 33416 3068 33468 3077
rect 35348 3136 35400 3188
rect 36636 3136 36688 3188
rect 37464 3179 37516 3188
rect 37464 3145 37473 3179
rect 37473 3145 37507 3179
rect 37507 3145 37516 3179
rect 37464 3136 37516 3145
rect 37556 3068 37608 3120
rect 5908 3000 5960 3052
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 11704 3043 11756 3052
rect 11704 3009 11713 3043
rect 11713 3009 11747 3043
rect 11747 3009 11756 3043
rect 11704 3000 11756 3009
rect 16212 3000 16264 3052
rect 18144 3043 18196 3052
rect 18144 3009 18153 3043
rect 18153 3009 18187 3043
rect 18187 3009 18196 3043
rect 18144 3000 18196 3009
rect 27804 3043 27856 3052
rect 27804 3009 27813 3043
rect 27813 3009 27847 3043
rect 27847 3009 27856 3043
rect 27804 3000 27856 3009
rect 33232 3043 33284 3052
rect 33232 3009 33241 3043
rect 33241 3009 33275 3043
rect 33275 3009 33284 3043
rect 33232 3000 33284 3009
rect 37648 3000 37700 3052
rect 3240 2932 3292 2984
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 12256 2975 12308 2984
rect 6460 2864 6512 2916
rect 12256 2941 12265 2975
rect 12265 2941 12299 2975
rect 12299 2941 12308 2975
rect 12256 2932 12308 2941
rect 18696 2975 18748 2984
rect 18696 2941 18705 2975
rect 18705 2941 18739 2975
rect 18739 2941 18748 2975
rect 18696 2932 18748 2941
rect 24492 2975 24544 2984
rect 24492 2941 24501 2975
rect 24501 2941 24535 2975
rect 24535 2941 24544 2975
rect 24492 2932 24544 2941
rect 28356 2975 28408 2984
rect 18788 2864 18840 2916
rect 28356 2941 28365 2975
rect 28365 2941 28399 2975
rect 28399 2941 28408 2975
rect 28356 2932 28408 2941
rect 35532 2932 35584 2984
rect 32588 2864 32640 2916
rect 5632 2796 5684 2848
rect 22192 2796 22244 2848
rect 32680 2796 32732 2848
rect 33692 2796 33744 2848
rect 35348 2796 35400 2848
rect 35992 2839 36044 2848
rect 35992 2805 36001 2839
rect 36001 2805 36035 2839
rect 36035 2805 36044 2839
rect 35992 2796 36044 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 21732 2592 21784 2644
rect 38108 2592 38160 2644
rect 4528 2524 4580 2576
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 1584 2499 1636 2508
rect 1584 2465 1593 2499
rect 1593 2465 1627 2499
rect 1627 2465 1636 2499
rect 1584 2456 1636 2465
rect 2780 2499 2832 2508
rect 2780 2465 2789 2499
rect 2789 2465 2823 2499
rect 2823 2465 2832 2499
rect 2780 2456 2832 2465
rect 5632 2499 5684 2508
rect 5632 2465 5641 2499
rect 5641 2465 5675 2499
rect 5675 2465 5684 2499
rect 5632 2456 5684 2465
rect 5816 2499 5868 2508
rect 5816 2465 5825 2499
rect 5825 2465 5859 2499
rect 5859 2465 5868 2499
rect 5816 2456 5868 2465
rect 6184 2456 6236 2508
rect 6552 2499 6604 2508
rect 6552 2465 6561 2499
rect 6561 2465 6595 2499
rect 6595 2465 6604 2499
rect 6552 2456 6604 2465
rect 9864 2524 9916 2576
rect 9312 2456 9364 2508
rect 9680 2499 9732 2508
rect 9680 2465 9689 2499
rect 9689 2465 9723 2499
rect 9723 2465 9732 2499
rect 9680 2456 9732 2465
rect 33692 2499 33744 2508
rect 33692 2465 33701 2499
rect 33701 2465 33735 2499
rect 33735 2465 33744 2499
rect 33692 2456 33744 2465
rect 37372 2524 37424 2576
rect 35992 2456 36044 2508
rect 21272 2388 21324 2440
rect 3884 2320 3936 2372
rect 35716 2320 35768 2372
rect 36728 2363 36780 2372
rect 36728 2329 36737 2363
rect 36737 2329 36771 2363
rect 36771 2329 36780 2363
rect 36728 2320 36780 2329
rect 37280 2252 37332 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect -10 49200 102 50000
rect 634 49200 746 50000
rect 1278 49200 1390 50000
rect 2566 49200 2678 50000
rect 2962 49736 3018 49745
rect 2962 49671 3018 49680
rect 32 46034 60 49200
rect 1398 47696 1454 47705
rect 1398 47631 1454 47640
rect 1412 47122 1440 47631
rect 1400 47116 1452 47122
rect 1400 47058 1452 47064
rect 2608 46646 2636 49200
rect 2872 47116 2924 47122
rect 2872 47058 2924 47064
rect 2596 46640 2648 46646
rect 2596 46582 2648 46588
rect 2780 46504 2832 46510
rect 2780 46446 2832 46452
rect 20 46028 72 46034
rect 20 45970 72 45976
rect 2792 45558 2820 46446
rect 2780 45552 2832 45558
rect 2780 45494 2832 45500
rect 1400 45416 1452 45422
rect 1400 45358 1452 45364
rect 1676 45416 1728 45422
rect 1676 45358 1728 45364
rect 1412 44985 1440 45358
rect 1398 44976 1454 44985
rect 1398 44911 1454 44920
rect 1584 43104 1636 43110
rect 1584 43046 1636 43052
rect 1596 42770 1624 43046
rect 1584 42764 1636 42770
rect 1584 42706 1636 42712
rect 1584 42628 1636 42634
rect 1584 42570 1636 42576
rect 1596 42362 1624 42570
rect 1584 42356 1636 42362
rect 1584 42298 1636 42304
rect 1400 41608 1452 41614
rect 1398 41576 1400 41585
rect 1452 41576 1454 41585
rect 1398 41511 1454 41520
rect 1584 40520 1636 40526
rect 1584 40462 1636 40468
rect 1596 40050 1624 40462
rect 1584 40044 1636 40050
rect 1584 39986 1636 39992
rect 1688 39030 1716 45358
rect 2884 45082 2912 47058
rect 2976 46510 3004 49671
rect 3210 49200 3322 50000
rect 3854 49200 3966 50000
rect 5142 49200 5254 50000
rect 5786 49200 5898 50000
rect 6430 49200 6542 50000
rect 7074 49314 7186 50000
rect 7074 49286 7512 49314
rect 7074 49200 7186 49286
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 3332 47184 3384 47190
rect 3332 47126 3384 47132
rect 3344 47025 3372 47126
rect 5184 47122 5212 49200
rect 4896 47116 4948 47122
rect 4896 47058 4948 47064
rect 5172 47116 5224 47122
rect 5172 47058 5224 47064
rect 3330 47016 3386 47025
rect 3056 46980 3108 46986
rect 3330 46951 3386 46960
rect 4620 46980 4672 46986
rect 3056 46922 3108 46928
rect 4620 46922 4672 46928
rect 2964 46504 3016 46510
rect 2964 46446 3016 46452
rect 3068 46170 3096 46922
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4632 46170 4660 46922
rect 4908 46170 4936 47058
rect 5448 46504 5500 46510
rect 5448 46446 5500 46452
rect 3056 46164 3108 46170
rect 3056 46106 3108 46112
rect 4620 46164 4672 46170
rect 4620 46106 4672 46112
rect 4896 46164 4948 46170
rect 4896 46106 4948 46112
rect 3240 45960 3292 45966
rect 3240 45902 3292 45908
rect 4804 45960 4856 45966
rect 4804 45902 4856 45908
rect 3056 45892 3108 45898
rect 3056 45834 3108 45840
rect 2964 45484 3016 45490
rect 2964 45426 3016 45432
rect 2976 45354 3004 45426
rect 2964 45348 3016 45354
rect 2964 45290 3016 45296
rect 2872 45076 2924 45082
rect 2872 45018 2924 45024
rect 2504 44872 2556 44878
rect 2504 44814 2556 44820
rect 2976 44826 3004 45290
rect 3068 45014 3096 45834
rect 3252 45490 3280 45902
rect 3240 45484 3292 45490
rect 3240 45426 3292 45432
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 3056 45008 3108 45014
rect 3056 44950 3108 44956
rect 2516 44742 2544 44814
rect 2976 44798 3096 44826
rect 2504 44736 2556 44742
rect 2504 44678 2556 44684
rect 2044 43104 2096 43110
rect 2044 43046 2096 43052
rect 2056 42226 2084 43046
rect 2044 42220 2096 42226
rect 2044 42162 2096 42168
rect 1768 39976 1820 39982
rect 1768 39918 1820 39924
rect 1780 39642 1808 39918
rect 1768 39636 1820 39642
rect 1768 39578 1820 39584
rect 2136 39432 2188 39438
rect 2136 39374 2188 39380
rect 1676 39024 1728 39030
rect 1676 38966 1728 38972
rect 1860 38888 1912 38894
rect 1860 38830 1912 38836
rect 1872 38554 1900 38830
rect 1860 38548 1912 38554
rect 1860 38490 1912 38496
rect 1400 36168 1452 36174
rect 1398 36136 1400 36145
rect 1452 36136 1454 36145
rect 1398 36071 1454 36080
rect 2148 30938 2176 39374
rect 2136 30932 2188 30938
rect 2136 30874 2188 30880
rect 1676 29640 1728 29646
rect 1676 29582 1728 29588
rect 1688 29170 1716 29582
rect 1676 29164 1728 29170
rect 1676 29106 1728 29112
rect 1860 29096 1912 29102
rect 1860 29038 1912 29044
rect 1872 28762 1900 29038
rect 1860 28756 1912 28762
rect 1860 28698 1912 28704
rect 2320 28552 2372 28558
rect 2320 28494 2372 28500
rect 1768 23112 1820 23118
rect 1768 23054 1820 23060
rect 1780 22642 1808 23054
rect 1952 22976 2004 22982
rect 1952 22918 2004 22924
rect 1964 22710 1992 22918
rect 1952 22704 2004 22710
rect 1952 22646 2004 22652
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1860 22092 1912 22098
rect 1860 22034 1912 22040
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1412 21146 1440 21966
rect 1872 21865 1900 22034
rect 2044 21956 2096 21962
rect 2044 21898 2096 21904
rect 1858 21856 1914 21865
rect 1858 21791 1914 21800
rect 2056 21690 2084 21898
rect 2044 21684 2096 21690
rect 2044 21626 2096 21632
rect 1400 21140 1452 21146
rect 1400 21082 1452 21088
rect 2332 20602 2360 28494
rect 2412 21548 2464 21554
rect 2412 21490 2464 21496
rect 2320 20596 2372 20602
rect 2320 20538 2372 20544
rect 1400 20256 1452 20262
rect 1400 20198 1452 20204
rect 1412 19922 1440 20198
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1860 19916 1912 19922
rect 1860 19858 1912 19864
rect 1872 19825 1900 19858
rect 1858 19816 1914 19825
rect 1858 19751 1914 19760
rect 1952 19780 2004 19786
rect 1952 19722 2004 19728
rect 1964 19514 1992 19722
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 2044 19372 2096 19378
rect 2044 19314 2096 19320
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1688 17746 1716 18022
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 2056 17218 2084 19314
rect 2136 17604 2188 17610
rect 2136 17546 2188 17552
rect 2148 17338 2176 17546
rect 2136 17332 2188 17338
rect 2136 17274 2188 17280
rect 2056 17190 2176 17218
rect 1400 16992 1452 16998
rect 1400 16934 1452 16940
rect 1412 16658 1440 16934
rect 1400 16652 1452 16658
rect 1400 16594 1452 16600
rect 1860 16652 1912 16658
rect 1860 16594 1912 16600
rect 1872 16425 1900 16594
rect 2044 16516 2096 16522
rect 2044 16458 2096 16464
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 2056 16250 2084 16458
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2148 16114 2176 17190
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 1398 15736 1454 15745
rect 1398 15671 1454 15680
rect 1412 15570 1440 15671
rect 1400 15564 1452 15570
rect 1400 15506 1452 15512
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1688 13938 1716 14350
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1872 13530 1900 13806
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1688 12850 1716 13262
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1860 12776 1912 12782
rect 1860 12718 1912 12724
rect 1872 12442 1900 12718
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 2148 11150 2176 16050
rect 2240 13326 2268 17138
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1596 10305 1624 10542
rect 1582 10296 1638 10305
rect 1582 10231 1638 10240
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1872 9586 1900 9998
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 2056 9654 2084 9862
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2056 8498 2084 8910
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2240 8566 2268 8774
rect 2228 8560 2280 8566
rect 2228 8502 2280 8508
rect 2044 8492 2096 8498
rect 2044 8434 2096 8440
rect 1400 8288 1452 8294
rect 1400 8230 1452 8236
rect 1412 7954 1440 8230
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 2228 7812 2280 7818
rect 2228 7754 2280 7760
rect 2240 7546 2268 7754
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 1400 7200 1452 7206
rect 1400 7142 1452 7148
rect 1412 6866 1440 7142
rect 1400 6860 1452 6866
rect 1400 6802 1452 6808
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 2056 6458 2084 6666
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 1400 5636 1452 5642
rect 1400 5578 1452 5584
rect 1412 5545 1440 5578
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 664 4004 716 4010
rect 664 3946 716 3952
rect 676 800 704 3946
rect 1412 2514 1440 4558
rect 1952 4072 2004 4078
rect 1952 4014 2004 4020
rect 1584 3392 1636 3398
rect 1584 3334 1636 3340
rect 1596 2514 1624 3334
rect 1964 3058 1992 4014
rect 2148 3534 2176 6258
rect 2332 5234 2360 14962
rect 2424 6322 2452 21490
rect 2516 10062 2544 44678
rect 2778 43616 2834 43625
rect 2778 43551 2834 43560
rect 2792 42770 2820 43551
rect 2780 42764 2832 42770
rect 2780 42706 2832 42712
rect 2962 42256 3018 42265
rect 2962 42191 3018 42200
rect 2976 42158 3004 42191
rect 2872 42152 2924 42158
rect 2872 42094 2924 42100
rect 2964 42152 3016 42158
rect 2964 42094 3016 42100
rect 2884 41818 2912 42094
rect 3068 41970 3096 44798
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 2976 41942 3096 41970
rect 2872 41812 2924 41818
rect 2872 41754 2924 41760
rect 2780 38888 2832 38894
rect 2872 38888 2924 38894
rect 2780 38830 2832 38836
rect 2870 38856 2872 38865
rect 2924 38856 2926 38865
rect 2792 38554 2820 38830
rect 2870 38791 2926 38800
rect 2780 38548 2832 38554
rect 2780 38490 2832 38496
rect 2778 29336 2834 29345
rect 2778 29271 2834 29280
rect 2792 29102 2820 29271
rect 2780 29096 2832 29102
rect 2780 29038 2832 29044
rect 2976 26234 3004 41942
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 3422 40896 3478 40905
rect 3422 40831 3478 40840
rect 3436 40118 3464 40831
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 3424 40112 3476 40118
rect 3424 40054 3476 40060
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4712 38344 4764 38350
rect 4712 38286 4764 38292
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 3330 37496 3386 37505
rect 4214 37488 4522 37508
rect 3330 37431 3386 37440
rect 3344 37330 3372 37431
rect 4724 37398 4752 38286
rect 4712 37392 4764 37398
rect 4712 37334 4764 37340
rect 3332 37324 3384 37330
rect 3332 37266 3384 37272
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 3240 36168 3292 36174
rect 3240 36110 3292 36116
rect 3056 36100 3108 36106
rect 3056 36042 3108 36048
rect 3068 35834 3096 36042
rect 3056 35828 3108 35834
rect 3056 35770 3108 35776
rect 3252 35630 3280 36110
rect 3240 35624 3292 35630
rect 3240 35566 3292 35572
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 2884 26206 3004 26234
rect 2780 22568 2832 22574
rect 2778 22536 2780 22545
rect 2832 22536 2834 22545
rect 2778 22471 2834 22480
rect 2778 17776 2834 17785
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13705 2820 13806
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2778 13016 2834 13025
rect 2778 12951 2834 12960
rect 2792 12782 2820 12951
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2778 9616 2834 9625
rect 2778 9551 2834 9560
rect 2792 9518 2820 9551
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2884 8974 2912 26206
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 3240 15904 3292 15910
rect 3240 15846 3292 15852
rect 3252 15570 3280 15846
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 3056 15428 3108 15434
rect 3056 15370 3108 15376
rect 3068 15162 3096 15370
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3252 10742 3280 11018
rect 3240 10736 3292 10742
rect 3240 10678 3292 10684
rect 3436 10674 3464 11086
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2778 8256 2834 8265
rect 2778 8191 2834 8200
rect 2792 7954 2820 8191
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2778 6896 2834 6905
rect 2778 6831 2780 6840
rect 2832 6831 2834 6840
rect 2780 6802 2832 6808
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2516 3738 2544 4014
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 2792 2145 2820 2450
rect 2778 2136 2834 2145
rect 2778 2071 2834 2080
rect 2884 1465 2912 8366
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3252 5778 3280 6054
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 3068 5370 3096 5578
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 3884 5160 3936 5166
rect 3884 5102 3936 5108
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 2976 4826 3004 5102
rect 3896 4826 3924 5102
rect 3988 4865 4016 5102
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 3974 4856 4030 4865
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 3884 4820 3936 4826
rect 4214 4848 4522 4868
rect 3974 4791 4030 4800
rect 3884 4762 3936 4768
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3988 4282 4016 4558
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 4080 4185 4108 4694
rect 4066 4176 4122 4185
rect 4724 4146 4752 37334
rect 4816 28490 4844 45902
rect 5460 43790 5488 46446
rect 5816 46368 5868 46374
rect 5816 46310 5868 46316
rect 6092 46368 6144 46374
rect 6092 46310 6144 46316
rect 5724 45892 5776 45898
rect 5724 45834 5776 45840
rect 5736 45626 5764 45834
rect 5724 45620 5776 45626
rect 5724 45562 5776 45568
rect 5828 45490 5856 46310
rect 6104 46034 6132 46310
rect 6472 46034 6500 49200
rect 7380 47116 7432 47122
rect 7380 47058 7432 47064
rect 6092 46028 6144 46034
rect 6092 45970 6144 45976
rect 6460 46028 6512 46034
rect 6460 45970 6512 45976
rect 6920 45552 6972 45558
rect 6920 45494 6972 45500
rect 5816 45484 5868 45490
rect 5816 45426 5868 45432
rect 6736 45416 6788 45422
rect 6736 45358 6788 45364
rect 6748 45082 6776 45358
rect 6736 45076 6788 45082
rect 6736 45018 6788 45024
rect 6932 44878 6960 45494
rect 7392 45082 7420 47058
rect 7484 45830 7512 49286
rect 8362 49200 8474 50000
rect 9006 49200 9118 50000
rect 9650 49200 9762 50000
rect 10938 49200 11050 50000
rect 11582 49200 11694 50000
rect 12226 49200 12338 50000
rect 12870 49200 12982 50000
rect 14158 49200 14270 50000
rect 14802 49200 14914 50000
rect 15446 49200 15558 50000
rect 16734 49200 16846 50000
rect 17378 49200 17490 50000
rect 18022 49200 18134 50000
rect 18666 49200 18778 50000
rect 19954 49200 20066 50000
rect 20598 49200 20710 50000
rect 21242 49200 21354 50000
rect 22530 49200 22642 50000
rect 23174 49200 23286 50000
rect 23818 49200 23930 50000
rect 24462 49200 24574 50000
rect 25750 49200 25862 50000
rect 26394 49200 26506 50000
rect 27038 49200 27150 50000
rect 28326 49200 28438 50000
rect 28970 49200 29082 50000
rect 29614 49200 29726 50000
rect 30258 49200 30370 50000
rect 31546 49200 31658 50000
rect 32190 49200 32302 50000
rect 32834 49200 32946 50000
rect 34122 49200 34234 50000
rect 34766 49200 34878 50000
rect 35410 49200 35522 50000
rect 36054 49450 36166 50000
rect 35912 49422 36166 49450
rect 8208 46980 8260 46986
rect 8208 46922 8260 46928
rect 8220 46714 8248 46922
rect 8208 46708 8260 46714
rect 8208 46650 8260 46656
rect 8404 46646 8432 49200
rect 8944 47048 8996 47054
rect 8944 46990 8996 46996
rect 8392 46640 8444 46646
rect 8392 46582 8444 46588
rect 8116 46572 8168 46578
rect 8116 46514 8168 46520
rect 8128 45966 8156 46514
rect 8208 46504 8260 46510
rect 8208 46446 8260 46452
rect 8220 46170 8248 46446
rect 8208 46164 8260 46170
rect 8208 46106 8260 46112
rect 8956 46034 8984 46990
rect 9048 46102 9076 49200
rect 9772 47048 9824 47054
rect 9772 46990 9824 46996
rect 9784 46578 9812 46990
rect 9772 46572 9824 46578
rect 9772 46514 9824 46520
rect 14924 46368 14976 46374
rect 14924 46310 14976 46316
rect 9036 46096 9088 46102
rect 9036 46038 9088 46044
rect 14936 46034 14964 46310
rect 15488 46034 15516 49200
rect 17420 47122 17448 49200
rect 18064 47410 18092 49200
rect 17972 47382 18092 47410
rect 17408 47116 17460 47122
rect 17408 47058 17460 47064
rect 16856 47048 16908 47054
rect 16856 46990 16908 46996
rect 16868 46578 16896 46990
rect 17040 46980 17092 46986
rect 17040 46922 17092 46928
rect 16856 46572 16908 46578
rect 16856 46514 16908 46520
rect 17052 46170 17080 46922
rect 17040 46164 17092 46170
rect 17040 46106 17092 46112
rect 8944 46028 8996 46034
rect 8944 45970 8996 45976
rect 14924 46028 14976 46034
rect 14924 45970 14976 45976
rect 15476 46028 15528 46034
rect 15476 45970 15528 45976
rect 8116 45960 8168 45966
rect 8036 45908 8116 45914
rect 8036 45902 8168 45908
rect 17408 45960 17460 45966
rect 17408 45902 17460 45908
rect 8036 45886 8156 45902
rect 8944 45892 8996 45898
rect 7472 45824 7524 45830
rect 7472 45766 7524 45772
rect 8036 45490 8064 45886
rect 8944 45834 8996 45840
rect 15200 45892 15252 45898
rect 15200 45834 15252 45840
rect 8116 45824 8168 45830
rect 8116 45766 8168 45772
rect 8024 45484 8076 45490
rect 8024 45426 8076 45432
rect 7380 45076 7432 45082
rect 7380 45018 7432 45024
rect 6920 44872 6972 44878
rect 6920 44814 6972 44820
rect 5448 43784 5500 43790
rect 5448 43726 5500 43732
rect 4804 28484 4856 28490
rect 4804 28426 4856 28432
rect 7840 27328 7892 27334
rect 7840 27270 7892 27276
rect 7852 26994 7880 27270
rect 8036 27130 8064 45426
rect 8128 45422 8156 45766
rect 8956 45626 8984 45834
rect 8944 45620 8996 45626
rect 8944 45562 8996 45568
rect 15212 45558 15240 45834
rect 15200 45552 15252 45558
rect 15200 45494 15252 45500
rect 8852 45484 8904 45490
rect 8852 45426 8904 45432
rect 15292 45484 15344 45490
rect 15292 45426 15344 45432
rect 8116 45416 8168 45422
rect 8116 45358 8168 45364
rect 8864 45082 8892 45426
rect 10048 45348 10100 45354
rect 10048 45290 10100 45296
rect 8852 45076 8904 45082
rect 8852 45018 8904 45024
rect 8208 44872 8260 44878
rect 8208 44814 8260 44820
rect 8024 27124 8076 27130
rect 8024 27066 8076 27072
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 7852 21554 7880 26930
rect 7840 21548 7892 21554
rect 7840 21490 7892 21496
rect 7852 20942 7880 21490
rect 8220 21010 8248 44814
rect 8864 41614 8892 45018
rect 9680 42220 9732 42226
rect 9680 42162 9732 42168
rect 9692 41614 9720 42162
rect 10060 41682 10088 45290
rect 10508 44736 10560 44742
rect 10508 44678 10560 44684
rect 10416 42152 10468 42158
rect 10416 42094 10468 42100
rect 10428 42022 10456 42094
rect 10416 42016 10468 42022
rect 10416 41958 10468 41964
rect 10048 41676 10100 41682
rect 10048 41618 10100 41624
rect 8852 41608 8904 41614
rect 8852 41550 8904 41556
rect 9680 41608 9732 41614
rect 9680 41550 9732 41556
rect 8392 41472 8444 41478
rect 8392 41414 8444 41420
rect 8404 41138 8432 41414
rect 8392 41132 8444 41138
rect 8392 41074 8444 41080
rect 8404 27470 8432 41074
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8864 26234 8892 41550
rect 9692 41206 9720 41550
rect 10060 41478 10088 41618
rect 10048 41472 10100 41478
rect 10048 41414 10100 41420
rect 9680 41200 9732 41206
rect 9680 41142 9732 41148
rect 9692 40526 9720 41142
rect 9680 40520 9732 40526
rect 9680 40462 9732 40468
rect 9692 40118 9720 40462
rect 9772 40180 9824 40186
rect 9772 40122 9824 40128
rect 9680 40112 9732 40118
rect 9680 40054 9732 40060
rect 9588 28484 9640 28490
rect 9588 28426 9640 28432
rect 9600 27674 9628 28426
rect 9588 27668 9640 27674
rect 9588 27610 9640 27616
rect 8772 26206 8892 26234
rect 8772 21486 8800 26206
rect 9600 23050 9628 27610
rect 9588 23044 9640 23050
rect 9588 22986 9640 22992
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8208 21004 8260 21010
rect 8208 20946 8260 20952
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7852 20534 7880 20878
rect 7840 20528 7892 20534
rect 7840 20470 7892 20476
rect 7852 19854 7880 20470
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 8116 19780 8168 19786
rect 8116 19722 8168 19728
rect 8128 18358 8156 19722
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 7012 7404 7064 7410
rect 7012 7346 7064 7352
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6380 4690 6408 4966
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 4066 4111 4122 4120
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 4816 3602 4844 3878
rect 5368 3670 5396 3878
rect 5356 3664 5408 3670
rect 5356 3606 5408 3612
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 2964 3460 3016 3466
rect 2964 3402 3016 3408
rect 2976 3058 3004 3402
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3160 3126 3188 3334
rect 3148 3120 3200 3126
rect 3148 3062 3200 3068
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 2870 1456 2926 1465
rect 2870 1391 2926 1400
rect 3252 800 3280 2926
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4528 2576 4580 2582
rect 4528 2518 4580 2524
rect 3884 2372 3936 2378
rect 3884 2314 3936 2320
rect 3896 800 3924 2314
rect 4540 800 4568 2518
rect 5184 800 5212 3538
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5644 2514 5672 2790
rect 5828 2514 5856 4490
rect 5920 3058 5948 4558
rect 5908 3052 5960 3058
rect 5908 2994 5960 3000
rect 6196 2514 6224 4626
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6644 3936 6696 3942
rect 6644 3878 6696 3884
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6472 800 6500 2858
rect 6564 2514 6592 3878
rect 6656 3505 6684 3878
rect 7024 3534 7052 7346
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7300 4146 7328 4490
rect 7392 4146 7420 18294
rect 8220 4622 8248 20946
rect 8772 11762 8800 21422
rect 9220 20392 9272 20398
rect 9220 20334 9272 20340
rect 9232 12434 9260 20334
rect 9232 12406 9444 12434
rect 9416 12238 9444 12406
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 8944 5024 8996 5030
rect 8944 4966 8996 4972
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8220 4162 8248 4558
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7380 4140 7432 4146
rect 8220 4134 8340 4162
rect 7380 4082 7432 4088
rect 7012 3528 7064 3534
rect 6642 3496 6698 3505
rect 7012 3470 7064 3476
rect 6642 3431 6698 3440
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 3126 6868 3334
rect 7116 3194 7144 4082
rect 7104 3188 7156 3194
rect 7104 3130 7156 3136
rect 8312 3126 8340 4134
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8680 3738 8708 4014
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8956 3058 8984 4966
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9140 3126 9168 3334
rect 9128 3120 9180 3126
rect 9128 3062 9180 3068
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 6552 2508 6604 2514
rect 6552 2450 6604 2456
rect 7116 800 7144 2926
rect 9324 2514 9352 4422
rect 9416 4078 9444 12174
rect 9496 4208 9548 4214
rect 9496 4150 9548 4156
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9508 4010 9536 4150
rect 9496 4004 9548 4010
rect 9496 3946 9548 3952
rect 9784 3534 9812 40122
rect 10428 12434 10456 41958
rect 10520 41274 10548 44678
rect 14464 42084 14516 42090
rect 14464 42026 14516 42032
rect 10508 41268 10560 41274
rect 10508 41210 10560 41216
rect 10968 40588 11020 40594
rect 10968 40530 11020 40536
rect 10980 37398 11008 40530
rect 14096 38752 14148 38758
rect 14096 38694 14148 38700
rect 14108 37874 14136 38694
rect 14096 37868 14148 37874
rect 14096 37810 14148 37816
rect 10968 37392 11020 37398
rect 10968 37334 11020 37340
rect 10980 31482 11008 37334
rect 14280 37324 14332 37330
rect 14280 37266 14332 37272
rect 14292 36854 14320 37266
rect 14280 36848 14332 36854
rect 14280 36790 14332 36796
rect 14372 36712 14424 36718
rect 14372 36654 14424 36660
rect 14384 36378 14412 36654
rect 14372 36372 14424 36378
rect 14372 36314 14424 36320
rect 14096 36168 14148 36174
rect 14096 36110 14148 36116
rect 14108 35698 14136 36110
rect 14096 35692 14148 35698
rect 14096 35634 14148 35640
rect 10968 31476 11020 31482
rect 10968 31418 11020 31424
rect 14108 29170 14136 35634
rect 14280 31136 14332 31142
rect 14280 31078 14332 31084
rect 14292 30734 14320 31078
rect 14280 30728 14332 30734
rect 14280 30670 14332 30676
rect 14188 29640 14240 29646
rect 14188 29582 14240 29588
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14200 28150 14228 29582
rect 14372 29504 14424 29510
rect 14372 29446 14424 29452
rect 14384 29170 14412 29446
rect 14372 29164 14424 29170
rect 14372 29106 14424 29112
rect 14188 28144 14240 28150
rect 14188 28086 14240 28092
rect 12900 28076 12952 28082
rect 12900 28018 12952 28024
rect 12912 27470 12940 28018
rect 14476 28014 14504 42026
rect 15304 40594 15332 45426
rect 16672 43716 16724 43722
rect 16672 43658 16724 43664
rect 16580 43240 16632 43246
rect 16580 43182 16632 43188
rect 16488 42560 16540 42566
rect 16488 42502 16540 42508
rect 16500 41614 16528 42502
rect 16592 42226 16620 43182
rect 16684 42770 16712 43658
rect 17224 43648 17276 43654
rect 17224 43590 17276 43596
rect 17236 43382 17264 43590
rect 17224 43376 17276 43382
rect 17224 43318 17276 43324
rect 16672 42764 16724 42770
rect 16672 42706 16724 42712
rect 16580 42220 16632 42226
rect 16580 42162 16632 42168
rect 16488 41608 16540 41614
rect 16488 41550 16540 41556
rect 16592 41546 16620 42162
rect 17420 41562 17448 45902
rect 17972 45422 18000 47382
rect 18708 46510 18736 49200
rect 19996 46918 20024 49200
rect 20812 47184 20864 47190
rect 20812 47126 20864 47132
rect 20168 47048 20220 47054
rect 20168 46990 20220 46996
rect 19984 46912 20036 46918
rect 19984 46854 20036 46860
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 18236 46504 18288 46510
rect 18236 46446 18288 46452
rect 18696 46504 18748 46510
rect 18696 46446 18748 46452
rect 18248 46170 18276 46446
rect 19432 46368 19484 46374
rect 19432 46310 19484 46316
rect 18236 46164 18288 46170
rect 18236 46106 18288 46112
rect 18052 45960 18104 45966
rect 18052 45902 18104 45908
rect 17960 45416 18012 45422
rect 17960 45358 18012 45364
rect 16580 41540 16632 41546
rect 16580 41482 16632 41488
rect 17420 41534 17724 41562
rect 18064 41546 18092 45902
rect 19340 45824 19392 45830
rect 19340 45766 19392 45772
rect 19352 45558 19380 45766
rect 19340 45552 19392 45558
rect 19340 45494 19392 45500
rect 19444 45422 19472 46310
rect 20180 46034 20208 46990
rect 20536 46572 20588 46578
rect 20536 46514 20588 46520
rect 20352 46368 20404 46374
rect 20352 46310 20404 46316
rect 20364 46034 20392 46310
rect 20168 46028 20220 46034
rect 20168 45970 20220 45976
rect 20352 46028 20404 46034
rect 20352 45970 20404 45976
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 20076 45484 20128 45490
rect 20076 45426 20128 45432
rect 19432 45416 19484 45422
rect 19432 45358 19484 45364
rect 19800 45416 19852 45422
rect 19800 45358 19852 45364
rect 19812 44946 19840 45358
rect 18144 44940 18196 44946
rect 18144 44882 18196 44888
rect 19800 44940 19852 44946
rect 19800 44882 19852 44888
rect 18156 44402 18184 44882
rect 19432 44872 19484 44878
rect 19432 44814 19484 44820
rect 18144 44396 18196 44402
rect 18144 44338 18196 44344
rect 19248 44396 19300 44402
rect 19248 44338 19300 44344
rect 19260 43994 19288 44338
rect 19444 44198 19472 44814
rect 19984 44736 20036 44742
rect 19984 44678 20036 44684
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19996 44402 20024 44678
rect 20088 44538 20116 45426
rect 20076 44532 20128 44538
rect 20076 44474 20128 44480
rect 19984 44396 20036 44402
rect 19984 44338 20036 44344
rect 19432 44192 19484 44198
rect 19432 44134 19484 44140
rect 20260 44192 20312 44198
rect 20260 44134 20312 44140
rect 19248 43988 19300 43994
rect 19248 43930 19300 43936
rect 19432 43784 19484 43790
rect 19432 43726 19484 43732
rect 19444 43450 19472 43726
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19432 43444 19484 43450
rect 19432 43386 19484 43392
rect 19984 43376 20036 43382
rect 19984 43318 20036 43324
rect 18236 43104 18288 43110
rect 18236 43046 18288 43052
rect 19248 43104 19300 43110
rect 19248 43046 19300 43052
rect 18248 41682 18276 43046
rect 18604 42696 18656 42702
rect 18604 42638 18656 42644
rect 18328 42560 18380 42566
rect 18328 42502 18380 42508
rect 18340 42226 18368 42502
rect 18328 42220 18380 42226
rect 18328 42162 18380 42168
rect 18616 41818 18644 42638
rect 19260 42566 19288 43046
rect 19996 42634 20024 43318
rect 20168 43308 20220 43314
rect 20168 43250 20220 43256
rect 20180 42838 20208 43250
rect 20272 43246 20300 44134
rect 20260 43240 20312 43246
rect 20260 43182 20312 43188
rect 20168 42832 20220 42838
rect 20168 42774 20220 42780
rect 19984 42628 20036 42634
rect 19984 42570 20036 42576
rect 19248 42560 19300 42566
rect 19248 42502 19300 42508
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19892 42016 19944 42022
rect 19996 42004 20024 42570
rect 20180 42362 20208 42774
rect 20272 42566 20300 43182
rect 20260 42560 20312 42566
rect 20260 42502 20312 42508
rect 20168 42356 20220 42362
rect 20168 42298 20220 42304
rect 19944 41976 20024 42004
rect 19892 41958 19944 41964
rect 18604 41812 18656 41818
rect 18604 41754 18656 41760
rect 20180 41682 20208 42298
rect 18236 41676 18288 41682
rect 18236 41618 18288 41624
rect 20168 41676 20220 41682
rect 20168 41618 20220 41624
rect 19432 41608 19484 41614
rect 19432 41550 19484 41556
rect 15292 40588 15344 40594
rect 15292 40530 15344 40536
rect 16764 40520 16816 40526
rect 16764 40462 16816 40468
rect 16672 40384 16724 40390
rect 16672 40326 16724 40332
rect 16684 40118 16712 40326
rect 16672 40112 16724 40118
rect 16672 40054 16724 40060
rect 16776 39642 16804 40462
rect 16764 39636 16816 39642
rect 16764 39578 16816 39584
rect 16856 39364 16908 39370
rect 16856 39306 16908 39312
rect 16868 38962 16896 39306
rect 16856 38956 16908 38962
rect 16856 38898 16908 38904
rect 16580 38752 16632 38758
rect 16580 38694 16632 38700
rect 16488 38344 16540 38350
rect 16488 38286 16540 38292
rect 15936 38276 15988 38282
rect 15936 38218 15988 38224
rect 15948 38010 15976 38218
rect 15936 38004 15988 38010
rect 15936 37946 15988 37952
rect 16500 37806 16528 38286
rect 16592 37874 16620 38694
rect 16580 37868 16632 37874
rect 16580 37810 16632 37816
rect 16764 37868 16816 37874
rect 16764 37810 16816 37816
rect 16488 37800 16540 37806
rect 16488 37742 16540 37748
rect 14648 37664 14700 37670
rect 14648 37606 14700 37612
rect 14660 37194 14688 37606
rect 16500 37262 16528 37742
rect 16776 37466 16804 37810
rect 16764 37460 16816 37466
rect 16764 37402 16816 37408
rect 16488 37256 16540 37262
rect 16488 37198 16540 37204
rect 14648 37188 14700 37194
rect 14648 37130 14700 37136
rect 16500 36786 16528 37198
rect 16856 37120 16908 37126
rect 16856 37062 16908 37068
rect 16488 36780 16540 36786
rect 16488 36722 16540 36728
rect 15752 36644 15804 36650
rect 15752 36586 15804 36592
rect 15568 35080 15620 35086
rect 15568 35022 15620 35028
rect 15580 34542 15608 35022
rect 15200 34536 15252 34542
rect 15200 34478 15252 34484
rect 15568 34536 15620 34542
rect 15568 34478 15620 34484
rect 15212 33930 15240 34478
rect 15108 33924 15160 33930
rect 15108 33866 15160 33872
rect 15200 33924 15252 33930
rect 15200 33866 15252 33872
rect 15120 33658 15148 33866
rect 15108 33652 15160 33658
rect 15108 33594 15160 33600
rect 15212 32502 15240 33866
rect 15384 33516 15436 33522
rect 15384 33458 15436 33464
rect 15396 33114 15424 33458
rect 15384 33108 15436 33114
rect 15384 33050 15436 33056
rect 15568 32904 15620 32910
rect 15568 32846 15620 32852
rect 15660 32904 15712 32910
rect 15660 32846 15712 32852
rect 15200 32496 15252 32502
rect 15200 32438 15252 32444
rect 14556 32428 14608 32434
rect 14556 32370 14608 32376
rect 14568 32026 14596 32370
rect 14556 32020 14608 32026
rect 14556 31962 14608 31968
rect 15580 31822 15608 32846
rect 15672 32570 15700 32846
rect 15660 32564 15712 32570
rect 15660 32506 15712 32512
rect 15568 31816 15620 31822
rect 15568 31758 15620 31764
rect 15580 31346 15608 31758
rect 15568 31340 15620 31346
rect 15568 31282 15620 31288
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 14936 29646 14964 30194
rect 15384 30184 15436 30190
rect 15384 30126 15436 30132
rect 14924 29640 14976 29646
rect 14924 29582 14976 29588
rect 14936 29170 14964 29582
rect 14924 29164 14976 29170
rect 14924 29106 14976 29112
rect 14648 28484 14700 28490
rect 14648 28426 14700 28432
rect 14464 28008 14516 28014
rect 14464 27950 14516 27956
rect 12900 27464 12952 27470
rect 12900 27406 12952 27412
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14200 19922 14228 23054
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14476 15026 14504 27950
rect 14660 27674 14688 28426
rect 14648 27668 14700 27674
rect 14648 27610 14700 27616
rect 14832 27532 14884 27538
rect 14832 27474 14884 27480
rect 14556 23044 14608 23050
rect 14556 22986 14608 22992
rect 14464 15020 14516 15026
rect 14464 14962 14516 14968
rect 10244 12406 10456 12434
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 9876 2582 9904 4558
rect 10244 3602 10272 12406
rect 14568 5302 14596 22986
rect 14556 5296 14608 5302
rect 14556 5238 14608 5244
rect 14844 4010 14872 27474
rect 14936 26994 14964 29106
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 15304 28082 15332 28494
rect 15292 28076 15344 28082
rect 15292 28018 15344 28024
rect 15304 27470 15332 28018
rect 15292 27464 15344 27470
rect 15292 27406 15344 27412
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 15200 26580 15252 26586
rect 15200 26522 15252 26528
rect 15212 21622 15240 26522
rect 15200 21616 15252 21622
rect 15200 21558 15252 21564
rect 15292 19780 15344 19786
rect 15292 19722 15344 19728
rect 15304 19310 15332 19722
rect 15292 19304 15344 19310
rect 15292 19246 15344 19252
rect 15396 17202 15424 30126
rect 15660 29708 15712 29714
rect 15660 29650 15712 29656
rect 15672 29617 15700 29650
rect 15658 29608 15714 29617
rect 15658 29543 15660 29552
rect 15712 29543 15714 29552
rect 15660 29514 15712 29520
rect 15672 29483 15700 29514
rect 15660 29096 15712 29102
rect 15658 29064 15660 29073
rect 15712 29064 15714 29073
rect 15658 28999 15714 29008
rect 15476 26920 15528 26926
rect 15476 26862 15528 26868
rect 15488 26586 15516 26862
rect 15476 26580 15528 26586
rect 15476 26522 15528 26528
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15672 24410 15700 24754
rect 15660 24404 15712 24410
rect 15660 24346 15712 24352
rect 15476 24200 15528 24206
rect 15476 24142 15528 24148
rect 15488 23254 15516 24142
rect 15568 23520 15620 23526
rect 15568 23462 15620 23468
rect 15660 23520 15712 23526
rect 15660 23462 15712 23468
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 15580 23118 15608 23462
rect 15672 23322 15700 23462
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 15764 22098 15792 36586
rect 15936 35012 15988 35018
rect 15936 34954 15988 34960
rect 15948 34746 15976 34954
rect 15936 34740 15988 34746
rect 15936 34682 15988 34688
rect 16500 34542 16528 36722
rect 16868 35894 16896 37062
rect 16776 35866 16896 35894
rect 17420 35894 17448 41534
rect 17696 41478 17724 41534
rect 18052 41540 18104 41546
rect 18052 41482 18104 41488
rect 19248 41540 19300 41546
rect 19248 41482 19300 41488
rect 17592 41472 17644 41478
rect 17592 41414 17644 41420
rect 17684 41472 17736 41478
rect 17684 41414 17736 41420
rect 17604 39506 17632 41414
rect 18696 40588 18748 40594
rect 18696 40530 18748 40536
rect 17868 40180 17920 40186
rect 17868 40122 17920 40128
rect 17592 39500 17644 39506
rect 17592 39442 17644 39448
rect 17604 38554 17632 39442
rect 17880 38894 17908 40122
rect 18144 40044 18196 40050
rect 18144 39986 18196 39992
rect 18156 39642 18184 39986
rect 18144 39636 18196 39642
rect 18144 39578 18196 39584
rect 18328 39432 18380 39438
rect 18328 39374 18380 39380
rect 18340 39098 18368 39374
rect 18708 39370 18736 40530
rect 18696 39364 18748 39370
rect 18696 39306 18748 39312
rect 18328 39092 18380 39098
rect 18328 39034 18380 39040
rect 18604 38956 18656 38962
rect 18604 38898 18656 38904
rect 17868 38888 17920 38894
rect 17868 38830 17920 38836
rect 17592 38548 17644 38554
rect 17592 38490 17644 38496
rect 17500 38208 17552 38214
rect 17500 38150 17552 38156
rect 17512 37942 17540 38150
rect 17500 37936 17552 37942
rect 17500 37878 17552 37884
rect 17512 37126 17540 37878
rect 17604 37194 17632 38490
rect 17880 38350 17908 38830
rect 18616 38418 18644 38898
rect 18144 38412 18196 38418
rect 18144 38354 18196 38360
rect 18604 38412 18656 38418
rect 18604 38354 18656 38360
rect 17868 38344 17920 38350
rect 17868 38286 17920 38292
rect 17776 38004 17828 38010
rect 17776 37946 17828 37952
rect 17788 37194 17816 37946
rect 17880 37398 17908 38286
rect 18156 38010 18184 38354
rect 18144 38004 18196 38010
rect 18144 37946 18196 37952
rect 18708 37874 18736 39306
rect 18696 37868 18748 37874
rect 18696 37810 18748 37816
rect 18512 37664 18564 37670
rect 18512 37606 18564 37612
rect 17868 37392 17920 37398
rect 17868 37334 17920 37340
rect 18524 37262 18552 37606
rect 18512 37256 18564 37262
rect 18512 37198 18564 37204
rect 17592 37188 17644 37194
rect 17592 37130 17644 37136
rect 17776 37188 17828 37194
rect 17776 37130 17828 37136
rect 17500 37120 17552 37126
rect 17500 37062 17552 37068
rect 17420 35866 17540 35894
rect 16672 34604 16724 34610
rect 16672 34546 16724 34552
rect 16488 34536 16540 34542
rect 16488 34478 16540 34484
rect 16684 34202 16712 34546
rect 16672 34196 16724 34202
rect 16672 34138 16724 34144
rect 16672 32564 16724 32570
rect 16672 32506 16724 32512
rect 16580 32292 16632 32298
rect 16580 32234 16632 32240
rect 16592 31770 16620 32234
rect 16684 31890 16712 32506
rect 16776 32434 16804 35866
rect 17408 35692 17460 35698
rect 17408 35634 17460 35640
rect 17224 35488 17276 35494
rect 17224 35430 17276 35436
rect 17236 34678 17264 35430
rect 17420 35290 17448 35634
rect 17408 35284 17460 35290
rect 17408 35226 17460 35232
rect 17224 34672 17276 34678
rect 17224 34614 17276 34620
rect 16856 33992 16908 33998
rect 16856 33934 16908 33940
rect 16868 33114 16896 33934
rect 16856 33108 16908 33114
rect 16856 33050 16908 33056
rect 16948 32836 17000 32842
rect 16948 32778 17000 32784
rect 16764 32428 16816 32434
rect 16764 32370 16816 32376
rect 16776 32026 16804 32370
rect 16960 32026 16988 32778
rect 17040 32428 17092 32434
rect 17040 32370 17092 32376
rect 16764 32020 16816 32026
rect 16764 31962 16816 31968
rect 16948 32020 17000 32026
rect 16948 31962 17000 31968
rect 16672 31884 16724 31890
rect 16672 31826 16724 31832
rect 16592 31754 16712 31770
rect 16592 31748 16724 31754
rect 16592 31742 16672 31748
rect 16672 31690 16724 31696
rect 16684 31278 16712 31690
rect 16776 31346 16804 31962
rect 17052 31958 17080 32370
rect 17040 31952 17092 31958
rect 17040 31894 17092 31900
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16672 31272 16724 31278
rect 16672 31214 16724 31220
rect 16684 30870 16712 31214
rect 17052 30870 17080 31894
rect 16672 30864 16724 30870
rect 16672 30806 16724 30812
rect 17040 30864 17092 30870
rect 17040 30806 17092 30812
rect 15936 28756 15988 28762
rect 15936 28698 15988 28704
rect 15948 28014 15976 28698
rect 17316 28484 17368 28490
rect 17316 28426 17368 28432
rect 16672 28416 16724 28422
rect 16672 28358 16724 28364
rect 15936 28008 15988 28014
rect 15934 27976 15936 27985
rect 15988 27976 15990 27985
rect 15934 27911 15990 27920
rect 16580 26444 16632 26450
rect 16580 26386 16632 26392
rect 16212 26376 16264 26382
rect 16212 26318 16264 26324
rect 15844 25968 15896 25974
rect 15842 25936 15844 25945
rect 15896 25936 15898 25945
rect 15842 25871 15898 25880
rect 16224 25702 16252 26318
rect 16592 25838 16620 26386
rect 16684 25906 16712 28358
rect 17328 28218 17356 28426
rect 17316 28212 17368 28218
rect 17316 28154 17368 28160
rect 17512 27538 17540 35866
rect 18708 35086 18736 37810
rect 19260 36310 19288 41482
rect 19444 41138 19472 41550
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19432 41132 19484 41138
rect 19432 41074 19484 41080
rect 19444 39930 19472 41074
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 20352 40180 20404 40186
rect 20352 40122 20404 40128
rect 20364 40050 20392 40122
rect 20352 40044 20404 40050
rect 20352 39986 20404 39992
rect 19524 39976 19576 39982
rect 19444 39924 19524 39930
rect 19444 39918 19576 39924
rect 19444 39902 19564 39918
rect 19444 39030 19472 39902
rect 20076 39296 20128 39302
rect 20076 39238 20128 39244
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19432 39024 19484 39030
rect 19432 38966 19484 38972
rect 19340 37664 19392 37670
rect 19340 37606 19392 37612
rect 19352 36786 19380 37606
rect 19444 37262 19472 38966
rect 19984 38956 20036 38962
rect 19984 38898 20036 38904
rect 19996 38554 20024 38898
rect 19984 38548 20036 38554
rect 19984 38490 20036 38496
rect 20088 38350 20116 39238
rect 20168 38956 20220 38962
rect 20168 38898 20220 38904
rect 20180 38486 20208 38898
rect 20364 38570 20392 39986
rect 20272 38554 20392 38570
rect 20272 38548 20404 38554
rect 20272 38542 20352 38548
rect 20168 38480 20220 38486
rect 20168 38422 20220 38428
rect 20076 38344 20128 38350
rect 20076 38286 20128 38292
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 20088 37874 20116 38286
rect 20272 38010 20300 38542
rect 20352 38490 20404 38496
rect 20352 38412 20404 38418
rect 20352 38354 20404 38360
rect 20260 38004 20312 38010
rect 20260 37946 20312 37952
rect 20364 37874 20392 38354
rect 20444 38276 20496 38282
rect 20444 38218 20496 38224
rect 20456 37942 20484 38218
rect 20444 37936 20496 37942
rect 20444 37878 20496 37884
rect 19524 37868 19576 37874
rect 19524 37810 19576 37816
rect 20076 37868 20128 37874
rect 20076 37810 20128 37816
rect 20352 37868 20404 37874
rect 20352 37810 20404 37816
rect 19432 37256 19484 37262
rect 19432 37198 19484 37204
rect 19536 37194 19564 37810
rect 20260 37256 20312 37262
rect 20260 37198 20312 37204
rect 19524 37188 19576 37194
rect 19524 37130 19576 37136
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 20272 36854 20300 37198
rect 20364 36922 20392 37810
rect 20456 37126 20484 37878
rect 20444 37120 20496 37126
rect 20444 37062 20496 37068
rect 20352 36916 20404 36922
rect 20352 36858 20404 36864
rect 20260 36848 20312 36854
rect 20260 36790 20312 36796
rect 19340 36780 19392 36786
rect 19340 36722 19392 36728
rect 20272 36378 20300 36790
rect 20444 36576 20496 36582
rect 20444 36518 20496 36524
rect 20260 36372 20312 36378
rect 20260 36314 20312 36320
rect 19248 36304 19300 36310
rect 19248 36246 19300 36252
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 20272 35894 20300 36314
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 20180 35866 20300 35894
rect 20180 35494 20208 35866
rect 20456 35766 20484 36518
rect 20444 35760 20496 35766
rect 20444 35702 20496 35708
rect 20168 35488 20220 35494
rect 20168 35430 20220 35436
rect 18328 35080 18380 35086
rect 18328 35022 18380 35028
rect 18696 35080 18748 35086
rect 18696 35022 18748 35028
rect 17868 35012 17920 35018
rect 17868 34954 17920 34960
rect 17880 34134 17908 34954
rect 18340 34746 18368 35022
rect 19248 34944 19300 34950
rect 19248 34886 19300 34892
rect 18328 34740 18380 34746
rect 18328 34682 18380 34688
rect 18144 34400 18196 34406
rect 18144 34342 18196 34348
rect 17868 34128 17920 34134
rect 17868 34070 17920 34076
rect 17880 33522 17908 34070
rect 18156 33998 18184 34342
rect 18340 33998 18368 34682
rect 19260 33998 19288 34886
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 19444 34202 19472 34546
rect 20180 34542 20208 35430
rect 20168 34536 20220 34542
rect 20168 34478 20220 34484
rect 19432 34196 19484 34202
rect 19432 34138 19484 34144
rect 20180 33998 20208 34478
rect 18144 33992 18196 33998
rect 18144 33934 18196 33940
rect 18328 33992 18380 33998
rect 18328 33934 18380 33940
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 20168 33992 20220 33998
rect 20168 33934 20220 33940
rect 18052 33856 18104 33862
rect 18052 33798 18104 33804
rect 17960 33652 18012 33658
rect 17960 33594 18012 33600
rect 17868 33516 17920 33522
rect 17868 33458 17920 33464
rect 17972 32910 18000 33594
rect 18064 33318 18092 33798
rect 18156 33454 18184 33934
rect 18340 33590 18368 33934
rect 18420 33856 18472 33862
rect 18420 33798 18472 33804
rect 20076 33856 20128 33862
rect 20076 33798 20128 33804
rect 18328 33584 18380 33590
rect 18328 33526 18380 33532
rect 18144 33448 18196 33454
rect 18144 33390 18196 33396
rect 18052 33312 18104 33318
rect 18052 33254 18104 33260
rect 17960 32904 18012 32910
rect 17960 32846 18012 32852
rect 18328 32428 18380 32434
rect 18328 32370 18380 32376
rect 18236 32224 18288 32230
rect 18236 32166 18288 32172
rect 18248 31822 18276 32166
rect 18340 32026 18368 32370
rect 18328 32020 18380 32026
rect 18328 31962 18380 31968
rect 18432 31890 18460 33798
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 18604 32972 18656 32978
rect 18604 32914 18656 32920
rect 18512 32768 18564 32774
rect 18512 32710 18564 32716
rect 18420 31884 18472 31890
rect 18420 31826 18472 31832
rect 18524 31822 18552 32710
rect 18616 32026 18644 32914
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 18604 32020 18656 32026
rect 18604 31962 18656 31968
rect 18236 31816 18288 31822
rect 18236 31758 18288 31764
rect 18512 31816 18564 31822
rect 18512 31758 18564 31764
rect 18420 31272 18472 31278
rect 18420 31214 18472 31220
rect 17684 31136 17736 31142
rect 17684 31078 17736 31084
rect 17696 30666 17724 31078
rect 18432 30734 18460 31214
rect 18052 30728 18104 30734
rect 18052 30670 18104 30676
rect 18420 30728 18472 30734
rect 18420 30670 18472 30676
rect 17684 30660 17736 30666
rect 17684 30602 17736 30608
rect 18064 29170 18092 30670
rect 18616 30258 18644 31962
rect 18696 31884 18748 31890
rect 18696 31826 18748 31832
rect 18708 31414 18736 31826
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 20088 31414 20116 33798
rect 20260 32224 20312 32230
rect 20260 32166 20312 32172
rect 20272 31822 20300 32166
rect 20260 31816 20312 31822
rect 20260 31758 20312 31764
rect 20548 31754 20576 46514
rect 20720 44872 20772 44878
rect 20720 44814 20772 44820
rect 20732 44470 20760 44814
rect 20720 44464 20772 44470
rect 20720 44406 20772 44412
rect 20824 42702 20852 47126
rect 21180 46572 21232 46578
rect 21180 46514 21232 46520
rect 21088 46368 21140 46374
rect 21088 46310 21140 46316
rect 20904 45280 20956 45286
rect 20904 45222 20956 45228
rect 20916 44402 20944 45222
rect 21100 44810 21128 46310
rect 21088 44804 21140 44810
rect 21088 44746 21140 44752
rect 21192 44538 21220 46514
rect 21284 46034 21312 49200
rect 22100 47048 22152 47054
rect 22100 46990 22152 46996
rect 22112 46578 22140 46990
rect 22572 46594 22600 49200
rect 24400 47048 24452 47054
rect 24400 46990 24452 46996
rect 22100 46572 22152 46578
rect 22572 46566 22692 46594
rect 24412 46578 24440 46990
rect 22100 46514 22152 46520
rect 22664 46510 22692 46566
rect 24400 46572 24452 46578
rect 24400 46514 24452 46520
rect 22560 46504 22612 46510
rect 22560 46446 22612 46452
rect 22652 46504 22704 46510
rect 22652 46446 22704 46452
rect 22572 46170 22600 46446
rect 24504 46442 24532 49200
rect 24584 46504 24636 46510
rect 24584 46446 24636 46452
rect 24492 46436 24544 46442
rect 24492 46378 24544 46384
rect 24596 46170 24624 46446
rect 26240 46368 26292 46374
rect 26240 46310 26292 46316
rect 22560 46164 22612 46170
rect 22560 46106 22612 46112
rect 24584 46164 24636 46170
rect 24584 46106 24636 46112
rect 26252 46034 26280 46310
rect 27080 46034 27108 49200
rect 27988 47048 28040 47054
rect 27988 46990 28040 46996
rect 28000 46578 28028 46990
rect 27988 46572 28040 46578
rect 27988 46514 28040 46520
rect 28368 46442 28396 49200
rect 29656 47138 29684 49200
rect 29656 47122 29776 47138
rect 29656 47116 29788 47122
rect 29656 47110 29736 47116
rect 29736 47058 29788 47064
rect 29552 47048 29604 47054
rect 29552 46990 29604 46996
rect 29276 46980 29328 46986
rect 29276 46922 29328 46928
rect 28632 46504 28684 46510
rect 28632 46446 28684 46452
rect 28356 46436 28408 46442
rect 28356 46378 28408 46384
rect 28644 46170 28672 46446
rect 28632 46164 28684 46170
rect 28632 46106 28684 46112
rect 21272 46028 21324 46034
rect 21272 45970 21324 45976
rect 26240 46028 26292 46034
rect 26240 45970 26292 45976
rect 27068 46028 27120 46034
rect 27068 45970 27120 45976
rect 22652 45960 22704 45966
rect 22652 45902 22704 45908
rect 23848 45960 23900 45966
rect 23848 45902 23900 45908
rect 28724 45960 28776 45966
rect 28724 45902 28776 45908
rect 22100 45484 22152 45490
rect 22100 45426 22152 45432
rect 22112 44742 22140 45426
rect 22192 45280 22244 45286
rect 22192 45222 22244 45228
rect 22100 44736 22152 44742
rect 22100 44678 22152 44684
rect 21180 44532 21232 44538
rect 21180 44474 21232 44480
rect 20904 44396 20956 44402
rect 20904 44338 20956 44344
rect 21456 44396 21508 44402
rect 21456 44338 21508 44344
rect 21468 43790 21496 44338
rect 22112 43858 22140 44678
rect 22100 43852 22152 43858
rect 22100 43794 22152 43800
rect 21456 43784 21508 43790
rect 21456 43726 21508 43732
rect 21180 43240 21232 43246
rect 21180 43182 21232 43188
rect 21192 42702 21220 43182
rect 21468 43178 21496 43726
rect 21456 43172 21508 43178
rect 21456 43114 21508 43120
rect 21272 43104 21324 43110
rect 21272 43046 21324 43052
rect 20812 42696 20864 42702
rect 20812 42638 20864 42644
rect 21180 42696 21232 42702
rect 21180 42638 21232 42644
rect 20996 42220 21048 42226
rect 20996 42162 21048 42168
rect 21008 41818 21036 42162
rect 20996 41812 21048 41818
rect 20996 41754 21048 41760
rect 20628 41472 20680 41478
rect 20628 41414 20680 41420
rect 20640 40934 20668 41414
rect 21192 41138 21220 42638
rect 21284 42634 21312 43046
rect 21468 42702 21496 43114
rect 22204 42702 22232 45222
rect 22376 44940 22428 44946
rect 22376 44882 22428 44888
rect 21456 42696 21508 42702
rect 21456 42638 21508 42644
rect 22192 42696 22244 42702
rect 22192 42638 22244 42644
rect 21272 42628 21324 42634
rect 21272 42570 21324 42576
rect 21272 42152 21324 42158
rect 21272 42094 21324 42100
rect 21284 41206 21312 42094
rect 21468 41546 21496 42638
rect 22284 42560 22336 42566
rect 22284 42502 22336 42508
rect 22296 42226 22324 42502
rect 22388 42226 22416 44882
rect 22664 42906 22692 45902
rect 23020 45484 23072 45490
rect 23020 45426 23072 45432
rect 22928 45348 22980 45354
rect 22928 45290 22980 45296
rect 22836 45280 22888 45286
rect 22836 45222 22888 45228
rect 22848 44742 22876 45222
rect 22940 44810 22968 45290
rect 23032 45014 23060 45426
rect 23020 45008 23072 45014
rect 23020 44950 23072 44956
rect 22928 44804 22980 44810
rect 22928 44746 22980 44752
rect 23032 44742 23060 44950
rect 23572 44872 23624 44878
rect 23572 44814 23624 44820
rect 23112 44804 23164 44810
rect 23112 44746 23164 44752
rect 22836 44736 22888 44742
rect 22836 44678 22888 44684
rect 23020 44736 23072 44742
rect 23020 44678 23072 44684
rect 23032 44538 23060 44678
rect 23020 44532 23072 44538
rect 23020 44474 23072 44480
rect 23124 43994 23152 44746
rect 23584 44402 23612 44814
rect 23664 44736 23716 44742
rect 23664 44678 23716 44684
rect 23676 44470 23704 44678
rect 23664 44464 23716 44470
rect 23664 44406 23716 44412
rect 23572 44396 23624 44402
rect 23572 44338 23624 44344
rect 23112 43988 23164 43994
rect 23112 43930 23164 43936
rect 22652 42900 22704 42906
rect 22652 42842 22704 42848
rect 22284 42220 22336 42226
rect 22284 42162 22336 42168
rect 22376 42220 22428 42226
rect 22376 42162 22428 42168
rect 22100 42016 22152 42022
rect 22100 41958 22152 41964
rect 21456 41540 21508 41546
rect 21456 41482 21508 41488
rect 21272 41200 21324 41206
rect 21272 41142 21324 41148
rect 21180 41132 21232 41138
rect 21180 41074 21232 41080
rect 20628 40928 20680 40934
rect 20628 40870 20680 40876
rect 21192 40526 21220 41074
rect 21284 40730 21312 41142
rect 21272 40724 21324 40730
rect 21272 40666 21324 40672
rect 21180 40520 21232 40526
rect 21180 40462 21232 40468
rect 21088 40452 21140 40458
rect 21088 40394 21140 40400
rect 20628 39976 20680 39982
rect 20628 39918 20680 39924
rect 20996 39976 21048 39982
rect 20996 39918 21048 39924
rect 20640 38418 20668 39918
rect 20812 39840 20864 39846
rect 20812 39782 20864 39788
rect 20824 38962 20852 39782
rect 20904 39364 20956 39370
rect 20904 39306 20956 39312
rect 20916 39098 20944 39306
rect 20904 39092 20956 39098
rect 20904 39034 20956 39040
rect 20812 38956 20864 38962
rect 20812 38898 20864 38904
rect 20904 38752 20956 38758
rect 20904 38694 20956 38700
rect 20628 38412 20680 38418
rect 20628 38354 20680 38360
rect 20720 37664 20772 37670
rect 20720 37606 20772 37612
rect 20628 37324 20680 37330
rect 20628 37266 20680 37272
rect 20640 36786 20668 37266
rect 20732 36854 20760 37606
rect 20916 36854 20944 38694
rect 20720 36848 20772 36854
rect 20720 36790 20772 36796
rect 20904 36848 20956 36854
rect 20904 36790 20956 36796
rect 20628 36780 20680 36786
rect 20628 36722 20680 36728
rect 20720 36712 20772 36718
rect 20720 36654 20772 36660
rect 20732 36038 20760 36654
rect 20904 36644 20956 36650
rect 20904 36586 20956 36592
rect 20720 36032 20772 36038
rect 20720 35974 20772 35980
rect 20628 32360 20680 32366
rect 20628 32302 20680 32308
rect 20640 31890 20668 32302
rect 20732 31958 20760 35974
rect 20916 35290 20944 36586
rect 20904 35284 20956 35290
rect 20904 35226 20956 35232
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20824 34746 20852 35022
rect 20812 34740 20864 34746
rect 20812 34682 20864 34688
rect 20916 33930 20944 35226
rect 21008 34592 21036 39918
rect 21100 36242 21128 40394
rect 21192 40050 21220 40462
rect 21180 40044 21232 40050
rect 21180 39986 21232 39992
rect 21284 39914 21312 40666
rect 22112 40458 22140 41958
rect 22100 40452 22152 40458
rect 22100 40394 22152 40400
rect 22664 40118 22692 42842
rect 23480 42764 23532 42770
rect 23480 42706 23532 42712
rect 23572 42764 23624 42770
rect 23572 42706 23624 42712
rect 22836 42560 22888 42566
rect 22836 42502 22888 42508
rect 22848 42226 22876 42502
rect 23296 42356 23348 42362
rect 23296 42298 23348 42304
rect 22836 42220 22888 42226
rect 22836 42162 22888 42168
rect 23308 42158 23336 42298
rect 22744 42152 22796 42158
rect 22744 42094 22796 42100
rect 23296 42152 23348 42158
rect 23296 42094 23348 42100
rect 22756 41818 22784 42094
rect 22744 41812 22796 41818
rect 22744 41754 22796 41760
rect 22756 41138 22784 41754
rect 22744 41132 22796 41138
rect 22744 41074 22796 41080
rect 22652 40112 22704 40118
rect 22652 40054 22704 40060
rect 21916 40044 21968 40050
rect 21916 39986 21968 39992
rect 21272 39908 21324 39914
rect 21272 39850 21324 39856
rect 21284 39506 21312 39850
rect 21272 39500 21324 39506
rect 21272 39442 21324 39448
rect 21284 38418 21312 39442
rect 21928 39438 21956 39986
rect 21916 39432 21968 39438
rect 21916 39374 21968 39380
rect 21824 39296 21876 39302
rect 21824 39238 21876 39244
rect 21732 38956 21784 38962
rect 21732 38898 21784 38904
rect 21272 38412 21324 38418
rect 21272 38354 21324 38360
rect 21180 38208 21232 38214
rect 21180 38150 21232 38156
rect 21192 37874 21220 38150
rect 21180 37868 21232 37874
rect 21180 37810 21232 37816
rect 21272 37664 21324 37670
rect 21272 37606 21324 37612
rect 21284 37194 21312 37606
rect 21272 37188 21324 37194
rect 21272 37130 21324 37136
rect 21640 36304 21692 36310
rect 21640 36246 21692 36252
rect 21088 36236 21140 36242
rect 21088 36178 21140 36184
rect 21272 35488 21324 35494
rect 21272 35430 21324 35436
rect 21284 34610 21312 35430
rect 21652 34610 21680 36246
rect 21088 34604 21140 34610
rect 21008 34564 21088 34592
rect 21088 34546 21140 34552
rect 21272 34604 21324 34610
rect 21640 34604 21692 34610
rect 21272 34546 21324 34552
rect 21468 34564 21640 34592
rect 20904 33924 20956 33930
rect 20904 33866 20956 33872
rect 21100 33590 21128 34546
rect 21088 33584 21140 33590
rect 21088 33526 21140 33532
rect 20996 33516 21048 33522
rect 20996 33458 21048 33464
rect 21008 32978 21036 33458
rect 20996 32972 21048 32978
rect 20996 32914 21048 32920
rect 21008 32434 21036 32914
rect 20996 32428 21048 32434
rect 20996 32370 21048 32376
rect 21284 31958 21312 34546
rect 20720 31952 20772 31958
rect 20720 31894 20772 31900
rect 21272 31952 21324 31958
rect 21272 31894 21324 31900
rect 20628 31884 20680 31890
rect 20628 31826 20680 31832
rect 20996 31884 21048 31890
rect 20996 31826 21048 31832
rect 20456 31726 20576 31754
rect 18696 31408 18748 31414
rect 18696 31350 18748 31356
rect 20076 31408 20128 31414
rect 20076 31350 20128 31356
rect 20088 30734 20116 31350
rect 20076 30728 20128 30734
rect 20076 30670 20128 30676
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 18604 30048 18656 30054
rect 18604 29990 18656 29996
rect 18616 29714 18644 29990
rect 18604 29708 18656 29714
rect 18604 29650 18656 29656
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 18236 29164 18288 29170
rect 18236 29106 18288 29112
rect 18064 28626 18092 29106
rect 18144 28960 18196 28966
rect 18144 28902 18196 28908
rect 18052 28620 18104 28626
rect 18052 28562 18104 28568
rect 18156 28558 18184 28902
rect 18248 28762 18276 29106
rect 18236 28756 18288 28762
rect 18236 28698 18288 28704
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 18512 28552 18564 28558
rect 18512 28494 18564 28500
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17604 28082 17632 28358
rect 17592 28076 17644 28082
rect 17592 28018 17644 28024
rect 17776 28076 17828 28082
rect 17776 28018 17828 28024
rect 17684 27940 17736 27946
rect 17684 27882 17736 27888
rect 17500 27532 17552 27538
rect 17500 27474 17552 27480
rect 17224 27464 17276 27470
rect 17224 27406 17276 27412
rect 16764 27396 16816 27402
rect 16764 27338 16816 27344
rect 16672 25900 16724 25906
rect 16672 25842 16724 25848
rect 16580 25832 16632 25838
rect 16580 25774 16632 25780
rect 16212 25696 16264 25702
rect 16212 25638 16264 25644
rect 15936 24608 15988 24614
rect 15936 24550 15988 24556
rect 15948 23866 15976 24550
rect 16028 24064 16080 24070
rect 16028 24006 16080 24012
rect 15936 23860 15988 23866
rect 15936 23802 15988 23808
rect 16040 23730 16068 24006
rect 15844 23724 15896 23730
rect 15844 23666 15896 23672
rect 16028 23724 16080 23730
rect 16028 23666 16080 23672
rect 15752 22092 15804 22098
rect 15752 22034 15804 22040
rect 15856 22030 15884 23666
rect 16120 22092 16172 22098
rect 16120 22034 16172 22040
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 15844 22024 15896 22030
rect 15844 21966 15896 21972
rect 15672 20466 15700 21966
rect 16132 21146 16160 22034
rect 16224 21622 16252 25638
rect 16592 25294 16620 25774
rect 16580 25288 16632 25294
rect 16580 25230 16632 25236
rect 16304 23792 16356 23798
rect 16304 23734 16356 23740
rect 16316 23118 16344 23734
rect 16304 23112 16356 23118
rect 16304 23054 16356 23060
rect 16488 23112 16540 23118
rect 16488 23054 16540 23060
rect 16500 22642 16528 23054
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16488 22092 16540 22098
rect 16488 22034 16540 22040
rect 16212 21616 16264 21622
rect 16212 21558 16264 21564
rect 16120 21140 16172 21146
rect 16120 21082 16172 21088
rect 16224 21010 16252 21558
rect 16500 21146 16528 22034
rect 16580 22024 16632 22030
rect 16580 21966 16632 21972
rect 16672 22024 16724 22030
rect 16672 21966 16724 21972
rect 16592 21690 16620 21966
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16212 21004 16264 21010
rect 16212 20946 16264 20952
rect 16500 20534 16528 21082
rect 16684 20942 16712 21966
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 15752 20528 15804 20534
rect 15752 20470 15804 20476
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15476 20256 15528 20262
rect 15476 20198 15528 20204
rect 15488 19378 15516 20198
rect 15764 20058 15792 20470
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 15856 20058 15884 20402
rect 15752 20052 15804 20058
rect 15752 19994 15804 20000
rect 15844 20052 15896 20058
rect 15844 19994 15896 20000
rect 15476 19372 15528 19378
rect 15476 19314 15528 19320
rect 15764 19310 15792 19994
rect 15856 19378 15884 19994
rect 16776 19514 16804 27338
rect 17236 27130 17264 27406
rect 17696 27384 17724 27882
rect 17788 27674 17816 28018
rect 17776 27668 17828 27674
rect 17776 27610 17828 27616
rect 18420 27532 18472 27538
rect 18420 27474 18472 27480
rect 18328 27464 18380 27470
rect 18328 27406 18380 27412
rect 17776 27396 17828 27402
rect 17696 27356 17776 27384
rect 17776 27338 17828 27344
rect 17788 27130 17816 27338
rect 17224 27124 17276 27130
rect 17224 27066 17276 27072
rect 17776 27124 17828 27130
rect 17776 27066 17828 27072
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 16868 26518 16896 26930
rect 18052 26920 18104 26926
rect 18052 26862 18104 26868
rect 16856 26512 16908 26518
rect 16856 26454 16908 26460
rect 18064 26382 18092 26862
rect 18340 26382 18368 27406
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 18328 26376 18380 26382
rect 18328 26318 18380 26324
rect 16856 26308 16908 26314
rect 16856 26250 16908 26256
rect 16868 24818 16896 26250
rect 16948 26240 17000 26246
rect 16948 26182 17000 26188
rect 16960 25906 16988 26182
rect 17052 26042 17080 26318
rect 17040 26036 17092 26042
rect 17040 25978 17092 25984
rect 16948 25900 17000 25906
rect 16948 25842 17000 25848
rect 16960 25430 16988 25842
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 16948 25424 17000 25430
rect 16948 25366 17000 25372
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16868 24206 16896 24754
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16960 24138 16988 25366
rect 17880 24818 17908 25774
rect 18064 25498 18092 26318
rect 18340 26042 18368 26318
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18052 25492 18104 25498
rect 18052 25434 18104 25440
rect 18340 25362 18368 25978
rect 18328 25356 18380 25362
rect 18328 25298 18380 25304
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 17868 24812 17920 24818
rect 17868 24754 17920 24760
rect 16948 24132 17000 24138
rect 16948 24074 17000 24080
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 17512 23322 17540 23666
rect 17880 23662 17908 24754
rect 18248 24206 18276 25230
rect 18236 24200 18288 24206
rect 18236 24142 18288 24148
rect 18248 23866 18276 24142
rect 18328 24064 18380 24070
rect 18328 24006 18380 24012
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 18340 23798 18368 24006
rect 18432 23866 18460 27474
rect 18524 27130 18552 28494
rect 18512 27124 18564 27130
rect 18512 27066 18564 27072
rect 18512 26308 18564 26314
rect 18512 26250 18564 26256
rect 18524 25498 18552 26250
rect 18512 25492 18564 25498
rect 18512 25434 18564 25440
rect 18420 23860 18472 23866
rect 18420 23802 18472 23808
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17500 23316 17552 23322
rect 17500 23258 17552 23264
rect 16948 22432 17000 22438
rect 16948 22374 17000 22380
rect 16960 22030 16988 22374
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 17512 21554 17540 23258
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17500 21548 17552 21554
rect 17500 21490 17552 21496
rect 17500 21412 17552 21418
rect 17500 21354 17552 21360
rect 17512 20874 17540 21354
rect 17500 20868 17552 20874
rect 17500 20810 17552 20816
rect 17512 20466 17540 20810
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 16856 20256 16908 20262
rect 16856 20198 16908 20204
rect 16868 19786 16896 20198
rect 17040 19848 17092 19854
rect 17040 19790 17092 19796
rect 16856 19780 16908 19786
rect 16856 19722 16908 19728
rect 16764 19508 16816 19514
rect 16764 19450 16816 19456
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 15752 19304 15804 19310
rect 15752 19246 15804 19252
rect 17052 18290 17080 19790
rect 17512 19786 17540 20402
rect 17880 19854 17908 22510
rect 18052 21684 18104 21690
rect 18052 21626 18104 21632
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17500 19780 17552 19786
rect 17500 19722 17552 19728
rect 17880 19446 17908 19790
rect 17972 19514 18000 20198
rect 18064 20058 18092 21626
rect 18616 20398 18644 29650
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19340 29006 19392 29012
rect 19340 28948 19392 28954
rect 19432 28960 19484 28966
rect 18696 28552 18748 28558
rect 18696 28494 18748 28500
rect 18708 28082 18736 28494
rect 18788 28484 18840 28490
rect 18788 28426 18840 28432
rect 18696 28076 18748 28082
rect 18696 28018 18748 28024
rect 18800 27402 18828 28426
rect 18788 27396 18840 27402
rect 18788 27338 18840 27344
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18800 26586 18828 26862
rect 18788 26580 18840 26586
rect 18788 26522 18840 26528
rect 19352 26450 19380 28948
rect 19432 28902 19484 28908
rect 19444 28626 19472 28902
rect 20456 28694 20484 31726
rect 20640 31346 20668 31826
rect 20628 31340 20680 31346
rect 20628 31282 20680 31288
rect 20640 30870 20668 31282
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20628 30864 20680 30870
rect 20628 30806 20680 30812
rect 20824 30734 20852 31214
rect 20812 30728 20864 30734
rect 20812 30670 20864 30676
rect 20904 30660 20956 30666
rect 20904 30602 20956 30608
rect 20916 30258 20944 30602
rect 20904 30252 20956 30258
rect 20824 30212 20904 30240
rect 20824 29646 20852 30212
rect 20904 30194 20956 30200
rect 21008 30190 21036 31826
rect 21284 31414 21312 31894
rect 21272 31408 21324 31414
rect 21272 31350 21324 31356
rect 21180 31136 21232 31142
rect 21180 31078 21232 31084
rect 21088 30592 21140 30598
rect 21088 30534 21140 30540
rect 21100 30394 21128 30534
rect 21088 30388 21140 30394
rect 21088 30330 21140 30336
rect 21100 30258 21128 30330
rect 21088 30252 21140 30258
rect 21088 30194 21140 30200
rect 20996 30184 21048 30190
rect 20996 30126 21048 30132
rect 20904 30116 20956 30122
rect 20904 30058 20956 30064
rect 20916 29646 20944 30058
rect 21008 29850 21036 30126
rect 20996 29844 21048 29850
rect 20996 29786 21048 29792
rect 21100 29646 21128 30194
rect 21192 30190 21220 31078
rect 21284 30802 21312 31350
rect 21272 30796 21324 30802
rect 21272 30738 21324 30744
rect 21180 30184 21232 30190
rect 21180 30126 21232 30132
rect 21364 30116 21416 30122
rect 21364 30058 21416 30064
rect 21272 30048 21324 30054
rect 21272 29990 21324 29996
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20904 29640 20956 29646
rect 20904 29582 20956 29588
rect 21088 29640 21140 29646
rect 21088 29582 21140 29588
rect 20628 29504 20680 29510
rect 20628 29446 20680 29452
rect 20444 28688 20496 28694
rect 20444 28630 20496 28636
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 19444 28082 19472 28562
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 20640 28150 20668 29446
rect 21284 28150 21312 29990
rect 21376 29782 21404 30058
rect 21364 29776 21416 29782
rect 21364 29718 21416 29724
rect 21468 28558 21496 34564
rect 21640 34546 21692 34552
rect 21548 30252 21600 30258
rect 21548 30194 21600 30200
rect 21560 29578 21588 30194
rect 21640 29708 21692 29714
rect 21640 29650 21692 29656
rect 21548 29572 21600 29578
rect 21548 29514 21600 29520
rect 21456 28552 21508 28558
rect 21456 28494 21508 28500
rect 20260 28144 20312 28150
rect 20260 28086 20312 28092
rect 20628 28144 20680 28150
rect 20628 28086 20680 28092
rect 21272 28144 21324 28150
rect 21272 28086 21324 28092
rect 19432 28076 19484 28082
rect 19432 28018 19484 28024
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 19432 27940 19484 27946
rect 19432 27882 19484 27888
rect 19444 27606 19472 27882
rect 20180 27674 20208 28018
rect 20168 27668 20220 27674
rect 20168 27610 20220 27616
rect 19432 27600 19484 27606
rect 19432 27542 19484 27548
rect 20076 27532 20128 27538
rect 20076 27474 20128 27480
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 19248 26308 19300 26314
rect 19248 26250 19300 26256
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19064 25696 19116 25702
rect 19064 25638 19116 25644
rect 19076 25362 19104 25638
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 19168 25158 19196 25842
rect 19156 25152 19208 25158
rect 19156 25094 19208 25100
rect 18696 23520 18748 23526
rect 18696 23462 18748 23468
rect 18708 22710 18736 23462
rect 18696 22704 18748 22710
rect 18696 22646 18748 22652
rect 19168 21486 19196 25094
rect 19260 24274 19288 26250
rect 19352 25702 19380 26386
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19340 25696 19392 25702
rect 19340 25638 19392 25644
rect 19352 25294 19380 25638
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19248 24268 19300 24274
rect 19248 24210 19300 24216
rect 19444 23730 19472 25774
rect 19996 25430 20024 27406
rect 20088 26994 20116 27474
rect 20272 27062 20300 28086
rect 20904 28076 20956 28082
rect 20904 28018 20956 28024
rect 20628 27464 20680 27470
rect 20628 27406 20680 27412
rect 20260 27056 20312 27062
rect 20260 26998 20312 27004
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 20088 26450 20116 26930
rect 20168 26852 20220 26858
rect 20168 26794 20220 26800
rect 20076 26444 20128 26450
rect 20076 26386 20128 26392
rect 19984 25424 20036 25430
rect 19984 25366 20036 25372
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 20180 24206 20208 26794
rect 20272 26450 20300 26998
rect 20640 26586 20668 27406
rect 20628 26580 20680 26586
rect 20628 26522 20680 26528
rect 20260 26444 20312 26450
rect 20260 26386 20312 26392
rect 20812 26308 20864 26314
rect 20812 26250 20864 26256
rect 20824 25922 20852 26250
rect 20916 26042 20944 28018
rect 21272 27872 21324 27878
rect 21272 27814 21324 27820
rect 21284 27538 21312 27814
rect 21272 27532 21324 27538
rect 21272 27474 21324 27480
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 21192 26382 21220 26726
rect 21088 26376 21140 26382
rect 21088 26318 21140 26324
rect 21180 26376 21232 26382
rect 21180 26318 21232 26324
rect 21100 26042 21128 26318
rect 21284 26194 21312 27474
rect 21468 27470 21496 28494
rect 21456 27464 21508 27470
rect 21456 27406 21508 27412
rect 21192 26166 21312 26194
rect 20904 26036 20956 26042
rect 20904 25978 20956 25984
rect 21088 26036 21140 26042
rect 21088 25978 21140 25984
rect 20824 25906 20944 25922
rect 20824 25900 20956 25906
rect 20824 25894 20904 25900
rect 20904 25842 20956 25848
rect 20812 25832 20864 25838
rect 20812 25774 20864 25780
rect 20824 25294 20852 25774
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20812 25288 20864 25294
rect 20812 25230 20864 25236
rect 20732 24818 20760 25230
rect 20720 24812 20772 24818
rect 20720 24754 20772 24760
rect 20536 24744 20588 24750
rect 20536 24686 20588 24692
rect 20444 24608 20496 24614
rect 20444 24550 20496 24556
rect 20456 24206 20484 24550
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 20444 24200 20496 24206
rect 20444 24142 20496 24148
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 20180 23798 20208 24142
rect 20168 23792 20220 23798
rect 20168 23734 20220 23740
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19444 23118 19472 23666
rect 19432 23112 19484 23118
rect 19432 23054 19484 23060
rect 19444 22778 19472 23054
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 20548 22574 20576 24686
rect 20536 22568 20588 22574
rect 20536 22510 20588 22516
rect 20548 22098 20576 22510
rect 20732 22166 20760 24754
rect 20824 22778 20852 25230
rect 20916 23730 20944 25842
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 21008 24410 21036 25230
rect 21088 24812 21140 24818
rect 21088 24754 21140 24760
rect 20996 24404 21048 24410
rect 20996 24346 21048 24352
rect 21100 23866 21128 24754
rect 21192 24410 21220 26166
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 21284 24818 21312 25978
rect 21272 24812 21324 24818
rect 21272 24754 21324 24760
rect 21284 24614 21312 24754
rect 21652 24750 21680 29650
rect 21640 24744 21692 24750
rect 21640 24686 21692 24692
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21180 24404 21232 24410
rect 21180 24346 21232 24352
rect 21088 23860 21140 23866
rect 21088 23802 21140 23808
rect 21192 23730 21220 24346
rect 21652 24274 21680 24686
rect 21640 24268 21692 24274
rect 21640 24210 21692 24216
rect 20904 23724 20956 23730
rect 20904 23666 20956 23672
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 20720 22160 20772 22166
rect 20720 22102 20772 22108
rect 20536 22092 20588 22098
rect 20536 22034 20588 22040
rect 20720 22024 20772 22030
rect 20916 22012 20944 22918
rect 21652 22642 21680 22918
rect 21640 22636 21692 22642
rect 21640 22578 21692 22584
rect 20772 21984 20944 22012
rect 20720 21966 20772 21972
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 20732 21690 20760 21966
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 19340 21616 19392 21622
rect 19340 21558 19392 21564
rect 19156 21480 19208 21486
rect 19352 21468 19380 21558
rect 19616 21548 19668 21554
rect 19536 21508 19616 21536
rect 19536 21468 19564 21508
rect 19616 21490 19668 21496
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19352 21440 19564 21468
rect 19156 21422 19208 21428
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18052 20052 18104 20058
rect 18052 19994 18104 20000
rect 18064 19666 18092 19994
rect 18616 19922 18644 20334
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 19444 19786 19472 21440
rect 19996 21146 20024 21490
rect 20352 21480 20404 21486
rect 20352 21422 20404 21428
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20364 20874 20392 21422
rect 20732 20942 20760 21626
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20352 20868 20404 20874
rect 20352 20810 20404 20816
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 20364 20058 20392 20810
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20168 19916 20220 19922
rect 20168 19858 20220 19864
rect 19432 19780 19484 19786
rect 19432 19722 19484 19728
rect 19248 19712 19300 19718
rect 18064 19638 18184 19666
rect 19248 19654 19300 19660
rect 17960 19508 18012 19514
rect 18012 19468 18092 19496
rect 17960 19450 18012 19456
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17972 18970 18000 19314
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 18064 18766 18092 19468
rect 18156 19310 18184 19638
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18156 18834 18184 19246
rect 19260 18970 19288 19654
rect 19444 19514 19472 19722
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19432 19508 19484 19514
rect 19432 19450 19484 19456
rect 19340 19372 19392 19378
rect 19340 19314 19392 19320
rect 19352 18970 19380 19314
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 18144 18828 18196 18834
rect 18144 18770 18196 18776
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17328 18290 17356 18566
rect 18156 18426 18184 18770
rect 19260 18766 19288 18906
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19352 18426 19380 18702
rect 18144 18420 18196 18426
rect 18144 18362 18196 18368
rect 19340 18420 19392 18426
rect 19340 18362 19392 18368
rect 19444 18290 19472 19450
rect 20088 18766 20116 19654
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 17316 18284 17368 18290
rect 17316 18226 17368 18232
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19996 18222 20024 18634
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 20180 18154 20208 19858
rect 20364 19854 20392 19994
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20364 19514 20392 19790
rect 20904 19712 20956 19718
rect 20904 19654 20956 19660
rect 20352 19508 20404 19514
rect 20352 19450 20404 19456
rect 20364 18834 20392 19450
rect 20352 18828 20404 18834
rect 20352 18770 20404 18776
rect 20916 18766 20944 19654
rect 20996 19372 21048 19378
rect 20996 19314 21048 19320
rect 21008 18970 21036 19314
rect 20996 18964 21048 18970
rect 20996 18906 21048 18912
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20168 18148 20220 18154
rect 20168 18090 20220 18096
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 15476 4684 15528 4690
rect 15476 4626 15528 4632
rect 15200 4616 15252 4622
rect 15200 4558 15252 4564
rect 13820 4004 13872 4010
rect 13820 3946 13872 3952
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 10428 3602 10456 3878
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 9864 2576 9916 2582
rect 9864 2518 9916 2524
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9680 2508 9732 2514
rect 9680 2450 9732 2456
rect 9692 800 9720 2450
rect 10980 800 11008 3538
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 11716 3058 11744 3334
rect 11900 3126 11928 3878
rect 13832 3194 13860 3946
rect 15212 3670 15240 4558
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15396 4282 15424 4490
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 15200 3664 15252 3670
rect 15200 3606 15252 3612
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12268 800 12296 2926
rect 15488 800 15516 4626
rect 15580 3534 15608 17138
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 15750 4312 15806 4321
rect 19574 4304 19882 4324
rect 15750 4247 15806 4256
rect 15764 4214 15792 4247
rect 15752 4208 15804 4214
rect 15752 4150 15804 4156
rect 20364 4146 20392 9998
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 15672 4049 15700 4082
rect 15658 4040 15714 4049
rect 15658 3975 15714 3984
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15672 3194 15700 3975
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 20168 3936 20220 3942
rect 20168 3878 20220 3884
rect 16764 3596 16816 3602
rect 16764 3538 16816 3544
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 16224 3058 16252 3470
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 16776 800 16804 3538
rect 18156 3058 18184 3878
rect 20180 3602 20208 3878
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 18788 3528 18840 3534
rect 18788 3470 18840 3476
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18340 3126 18368 3334
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 18144 3052 18196 3058
rect 18144 2994 18196 3000
rect 18696 2984 18748 2990
rect 18696 2926 18748 2932
rect 18708 800 18736 2926
rect 18800 2922 18828 3470
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 18788 2916 18840 2922
rect 18788 2858 18840 2864
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 20640 800 20668 3538
rect 21744 2650 21772 38898
rect 21836 38894 21864 39238
rect 21824 38888 21876 38894
rect 21824 38830 21876 38836
rect 23020 38276 23072 38282
rect 23020 38218 23072 38224
rect 23032 37466 23060 38218
rect 23112 37868 23164 37874
rect 23112 37810 23164 37816
rect 23124 37466 23152 37810
rect 23020 37460 23072 37466
rect 23020 37402 23072 37408
rect 23112 37460 23164 37466
rect 23112 37402 23164 37408
rect 22836 37324 22888 37330
rect 22836 37266 22888 37272
rect 22376 37256 22428 37262
rect 22376 37198 22428 37204
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 22388 36310 22416 37198
rect 22480 36922 22508 37198
rect 22468 36916 22520 36922
rect 22468 36858 22520 36864
rect 22376 36304 22428 36310
rect 22376 36246 22428 36252
rect 21824 36168 21876 36174
rect 21824 36110 21876 36116
rect 21836 33386 21864 36110
rect 22744 35080 22796 35086
rect 22744 35022 22796 35028
rect 22560 34944 22612 34950
rect 22560 34886 22612 34892
rect 22572 34746 22600 34886
rect 22560 34740 22612 34746
rect 22560 34682 22612 34688
rect 22756 34610 22784 35022
rect 22848 34678 22876 37266
rect 23112 35692 23164 35698
rect 23112 35634 23164 35640
rect 23124 35018 23152 35634
rect 23112 35012 23164 35018
rect 23112 34954 23164 34960
rect 22836 34672 22888 34678
rect 22836 34614 22888 34620
rect 22744 34604 22796 34610
rect 22744 34546 22796 34552
rect 22836 34536 22888 34542
rect 22836 34478 22888 34484
rect 22848 33402 22876 34478
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 23032 33522 23060 33934
rect 23020 33516 23072 33522
rect 23020 33458 23072 33464
rect 21824 33380 21876 33386
rect 21824 33322 21876 33328
rect 22756 33374 22876 33402
rect 22008 33312 22060 33318
rect 22008 33254 22060 33260
rect 22020 32026 22048 33254
rect 22008 32020 22060 32026
rect 22008 31962 22060 31968
rect 22756 31958 22784 33374
rect 22836 33312 22888 33318
rect 22836 33254 22888 33260
rect 22744 31952 22796 31958
rect 22744 31894 22796 31900
rect 21824 31340 21876 31346
rect 21824 31282 21876 31288
rect 21836 30734 21864 31282
rect 22468 31272 22520 31278
rect 22468 31214 22520 31220
rect 21824 30728 21876 30734
rect 21824 30670 21876 30676
rect 21916 30592 21968 30598
rect 21916 30534 21968 30540
rect 21928 30258 21956 30534
rect 22008 30388 22060 30394
rect 22008 30330 22060 30336
rect 22020 30274 22048 30330
rect 22020 30258 22140 30274
rect 21916 30252 21968 30258
rect 21916 30194 21968 30200
rect 22020 30252 22152 30258
rect 22020 30246 22100 30252
rect 21824 30048 21876 30054
rect 21824 29990 21876 29996
rect 21836 26994 21864 29990
rect 22020 29646 22048 30246
rect 22100 30194 22152 30200
rect 22376 30252 22428 30258
rect 22376 30194 22428 30200
rect 22192 30184 22244 30190
rect 22192 30126 22244 30132
rect 22204 29714 22232 30126
rect 22388 29782 22416 30194
rect 22376 29776 22428 29782
rect 22376 29718 22428 29724
rect 22192 29708 22244 29714
rect 22192 29650 22244 29656
rect 22008 29640 22060 29646
rect 22008 29582 22060 29588
rect 22480 29170 22508 31214
rect 22848 30734 22876 33254
rect 23032 32502 23060 33458
rect 23112 33380 23164 33386
rect 23112 33322 23164 33328
rect 23020 32496 23072 32502
rect 23020 32438 23072 32444
rect 23020 31952 23072 31958
rect 23020 31894 23072 31900
rect 23032 31414 23060 31894
rect 23020 31408 23072 31414
rect 23020 31350 23072 31356
rect 22836 30728 22888 30734
rect 22836 30670 22888 30676
rect 22836 29776 22888 29782
rect 22836 29718 22888 29724
rect 22468 29164 22520 29170
rect 22468 29106 22520 29112
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 22480 28626 22508 29106
rect 22756 28762 22784 29106
rect 22848 28966 22876 29718
rect 23124 29646 23152 33322
rect 23204 32428 23256 32434
rect 23204 32370 23256 32376
rect 23216 32026 23244 32370
rect 23204 32020 23256 32026
rect 23204 31962 23256 31968
rect 23308 30598 23336 42094
rect 23492 41682 23520 42706
rect 23480 41676 23532 41682
rect 23480 41618 23532 41624
rect 23584 41528 23612 42706
rect 23756 42560 23808 42566
rect 23756 42502 23808 42508
rect 23768 42226 23796 42502
rect 23756 42220 23808 42226
rect 23756 42162 23808 42168
rect 23860 42090 23888 45902
rect 26424 45892 26476 45898
rect 26424 45834 26476 45840
rect 26436 45626 26464 45834
rect 26424 45620 26476 45626
rect 26424 45562 26476 45568
rect 24768 45484 24820 45490
rect 24768 45426 24820 45432
rect 24952 45484 25004 45490
rect 24952 45426 25004 45432
rect 27160 45484 27212 45490
rect 27160 45426 27212 45432
rect 24780 44946 24808 45426
rect 24768 44940 24820 44946
rect 24768 44882 24820 44888
rect 24780 44402 24808 44882
rect 24964 44810 24992 45426
rect 26884 45280 26936 45286
rect 26884 45222 26936 45228
rect 26056 44872 26108 44878
rect 26056 44814 26108 44820
rect 24952 44804 25004 44810
rect 24952 44746 25004 44752
rect 25780 44804 25832 44810
rect 25780 44746 25832 44752
rect 23940 44396 23992 44402
rect 23940 44338 23992 44344
rect 24768 44396 24820 44402
rect 24768 44338 24820 44344
rect 23952 43314 23980 44338
rect 25792 43994 25820 44746
rect 26068 44402 26096 44814
rect 26056 44396 26108 44402
rect 26056 44338 26108 44344
rect 25964 44192 26016 44198
rect 25964 44134 26016 44140
rect 25780 43988 25832 43994
rect 25780 43930 25832 43936
rect 25976 43790 26004 44134
rect 26068 43858 26096 44338
rect 26240 44328 26292 44334
rect 26240 44270 26292 44276
rect 26056 43852 26108 43858
rect 26056 43794 26108 43800
rect 25780 43784 25832 43790
rect 25780 43726 25832 43732
rect 25964 43784 26016 43790
rect 25964 43726 26016 43732
rect 25136 43648 25188 43654
rect 25136 43590 25188 43596
rect 23940 43308 23992 43314
rect 23940 43250 23992 43256
rect 24032 43308 24084 43314
rect 24032 43250 24084 43256
rect 23952 42770 23980 43250
rect 23940 42764 23992 42770
rect 23940 42706 23992 42712
rect 23940 42628 23992 42634
rect 23940 42570 23992 42576
rect 23848 42084 23900 42090
rect 23848 42026 23900 42032
rect 23848 41676 23900 41682
rect 23848 41618 23900 41624
rect 23664 41608 23716 41614
rect 23664 41550 23716 41556
rect 23492 41500 23612 41528
rect 23492 41426 23520 41500
rect 23400 41398 23520 41426
rect 23400 41206 23428 41398
rect 23388 41200 23440 41206
rect 23388 41142 23440 41148
rect 23676 40730 23704 41550
rect 23664 40724 23716 40730
rect 23664 40666 23716 40672
rect 23664 40520 23716 40526
rect 23664 40462 23716 40468
rect 23676 40186 23704 40462
rect 23664 40180 23716 40186
rect 23664 40122 23716 40128
rect 23676 39982 23704 40122
rect 23664 39976 23716 39982
rect 23664 39918 23716 39924
rect 23572 37664 23624 37670
rect 23572 37606 23624 37612
rect 23664 37664 23716 37670
rect 23664 37606 23716 37612
rect 23584 37262 23612 37606
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 23480 37120 23532 37126
rect 23480 37062 23532 37068
rect 23492 36922 23520 37062
rect 23480 36916 23532 36922
rect 23480 36858 23532 36864
rect 23388 36848 23440 36854
rect 23388 36790 23440 36796
rect 23400 36582 23428 36790
rect 23584 36786 23612 37198
rect 23572 36780 23624 36786
rect 23572 36722 23624 36728
rect 23388 36576 23440 36582
rect 23388 36518 23440 36524
rect 23400 35222 23428 36518
rect 23676 35766 23704 37606
rect 23756 37188 23808 37194
rect 23756 37130 23808 37136
rect 23768 36786 23796 37130
rect 23756 36780 23808 36786
rect 23756 36722 23808 36728
rect 23664 35760 23716 35766
rect 23584 35720 23664 35748
rect 23388 35216 23440 35222
rect 23584 35193 23612 35720
rect 23664 35702 23716 35708
rect 23768 35578 23796 36722
rect 23860 36174 23888 41618
rect 23952 41414 23980 42570
rect 24044 42362 24072 43250
rect 25148 42702 25176 43590
rect 25792 43450 25820 43726
rect 25780 43444 25832 43450
rect 25780 43386 25832 43392
rect 26068 43382 26096 43794
rect 26056 43376 26108 43382
rect 26056 43318 26108 43324
rect 26252 43178 26280 44270
rect 26896 43790 26924 45222
rect 26976 44736 27028 44742
rect 26976 44678 27028 44684
rect 26988 44402 27016 44678
rect 27172 44538 27200 45426
rect 28356 45416 28408 45422
rect 28356 45358 28408 45364
rect 27344 45008 27396 45014
rect 27344 44950 27396 44956
rect 27160 44532 27212 44538
rect 27160 44474 27212 44480
rect 26976 44396 27028 44402
rect 26976 44338 27028 44344
rect 26884 43784 26936 43790
rect 26884 43726 26936 43732
rect 26896 43450 26924 43726
rect 27356 43450 27384 44950
rect 27804 44396 27856 44402
rect 27804 44338 27856 44344
rect 27816 43994 27844 44338
rect 27988 44192 28040 44198
rect 27988 44134 28040 44140
rect 27804 43988 27856 43994
rect 27804 43930 27856 43936
rect 27620 43784 27672 43790
rect 27620 43726 27672 43732
rect 26884 43444 26936 43450
rect 26884 43386 26936 43392
rect 27344 43444 27396 43450
rect 27344 43386 27396 43392
rect 26240 43172 26292 43178
rect 26240 43114 26292 43120
rect 26252 42906 26280 43114
rect 26240 42900 26292 42906
rect 26240 42842 26292 42848
rect 26896 42770 26924 43386
rect 27068 43308 27120 43314
rect 27068 43250 27120 43256
rect 26976 43172 27028 43178
rect 26976 43114 27028 43120
rect 26884 42764 26936 42770
rect 26884 42706 26936 42712
rect 26988 42702 27016 43114
rect 27080 42906 27108 43250
rect 27160 43104 27212 43110
rect 27160 43046 27212 43052
rect 27068 42900 27120 42906
rect 27068 42842 27120 42848
rect 25136 42696 25188 42702
rect 25136 42638 25188 42644
rect 26976 42696 27028 42702
rect 26976 42638 27028 42644
rect 24032 42356 24084 42362
rect 24032 42298 24084 42304
rect 27172 42226 27200 43046
rect 27356 42702 27384 43386
rect 27344 42696 27396 42702
rect 27344 42638 27396 42644
rect 27160 42220 27212 42226
rect 27160 42162 27212 42168
rect 26976 42016 27028 42022
rect 26976 41958 27028 41964
rect 26988 41614 27016 41958
rect 27632 41614 27660 43726
rect 28000 43722 28028 44134
rect 28368 43790 28396 45358
rect 28356 43784 28408 43790
rect 28356 43726 28408 43732
rect 27988 43716 28040 43722
rect 27988 43658 28040 43664
rect 27712 42560 27764 42566
rect 27712 42502 27764 42508
rect 27804 42560 27856 42566
rect 27804 42502 27856 42508
rect 27724 42294 27752 42502
rect 27816 42362 27844 42502
rect 27804 42356 27856 42362
rect 27804 42298 27856 42304
rect 27712 42288 27764 42294
rect 27712 42230 27764 42236
rect 27712 42152 27764 42158
rect 27712 42094 27764 42100
rect 26976 41608 27028 41614
rect 26976 41550 27028 41556
rect 27620 41608 27672 41614
rect 27620 41550 27672 41556
rect 26148 41472 26200 41478
rect 26148 41414 26200 41420
rect 23952 41386 24072 41414
rect 23940 38752 23992 38758
rect 23940 38694 23992 38700
rect 23952 37874 23980 38694
rect 23940 37868 23992 37874
rect 23940 37810 23992 37816
rect 23848 36168 23900 36174
rect 23848 36110 23900 36116
rect 24044 35834 24072 41386
rect 25228 41132 25280 41138
rect 25228 41074 25280 41080
rect 24860 40996 24912 41002
rect 24860 40938 24912 40944
rect 24872 40594 24900 40938
rect 25136 40928 25188 40934
rect 25136 40870 25188 40876
rect 24860 40588 24912 40594
rect 24860 40530 24912 40536
rect 24872 40050 24900 40530
rect 24952 40452 25004 40458
rect 24952 40394 25004 40400
rect 24860 40044 24912 40050
rect 24860 39986 24912 39992
rect 24964 39914 24992 40394
rect 24952 39908 25004 39914
rect 24952 39850 25004 39856
rect 24676 39840 24728 39846
rect 24676 39782 24728 39788
rect 24688 39438 24716 39782
rect 25044 39636 25096 39642
rect 25044 39578 25096 39584
rect 24676 39432 24728 39438
rect 24676 39374 24728 39380
rect 24688 38962 24716 39374
rect 25056 38962 25084 39578
rect 25148 39438 25176 40870
rect 25240 40458 25268 41074
rect 26056 40724 26108 40730
rect 26056 40666 26108 40672
rect 25872 40656 25924 40662
rect 25872 40598 25924 40604
rect 25228 40452 25280 40458
rect 25228 40394 25280 40400
rect 25596 40384 25648 40390
rect 25596 40326 25648 40332
rect 25780 40384 25832 40390
rect 25780 40326 25832 40332
rect 25608 39642 25636 40326
rect 25792 40050 25820 40326
rect 25884 40050 25912 40598
rect 25780 40044 25832 40050
rect 25780 39986 25832 39992
rect 25872 40044 25924 40050
rect 25872 39986 25924 39992
rect 25780 39840 25832 39846
rect 25780 39782 25832 39788
rect 25596 39636 25648 39642
rect 25596 39578 25648 39584
rect 25792 39506 25820 39782
rect 25780 39500 25832 39506
rect 25780 39442 25832 39448
rect 25136 39432 25188 39438
rect 25136 39374 25188 39380
rect 24676 38956 24728 38962
rect 24676 38898 24728 38904
rect 25044 38956 25096 38962
rect 25044 38898 25096 38904
rect 24688 38350 24716 38898
rect 25148 38826 25176 39374
rect 25320 39296 25372 39302
rect 25320 39238 25372 39244
rect 25228 38888 25280 38894
rect 25228 38830 25280 38836
rect 25136 38820 25188 38826
rect 25136 38762 25188 38768
rect 24860 38480 24912 38486
rect 24860 38422 24912 38428
rect 24872 38350 24900 38422
rect 25240 38418 25268 38830
rect 25228 38412 25280 38418
rect 25228 38354 25280 38360
rect 24676 38344 24728 38350
rect 24676 38286 24728 38292
rect 24860 38344 24912 38350
rect 24860 38286 24912 38292
rect 24216 38208 24268 38214
rect 24216 38150 24268 38156
rect 24860 38208 24912 38214
rect 24860 38150 24912 38156
rect 24228 37874 24256 38150
rect 24872 37942 24900 38150
rect 25332 37942 25360 39238
rect 25792 38962 25820 39442
rect 26068 38962 26096 40666
rect 26160 40662 26188 41414
rect 27724 41274 27752 42094
rect 28632 41608 28684 41614
rect 28632 41550 28684 41556
rect 26884 41268 26936 41274
rect 26884 41210 26936 41216
rect 27712 41268 27764 41274
rect 27712 41210 27764 41216
rect 26896 40934 26924 41210
rect 26976 41132 27028 41138
rect 26976 41074 27028 41080
rect 26884 40928 26936 40934
rect 26884 40870 26936 40876
rect 26148 40656 26200 40662
rect 26148 40598 26200 40604
rect 26988 40186 27016 41074
rect 27724 40526 27752 41210
rect 28644 41070 28672 41550
rect 27988 41064 28040 41070
rect 27988 41006 28040 41012
rect 28632 41064 28684 41070
rect 28632 41006 28684 41012
rect 28000 40526 28028 41006
rect 27712 40520 27764 40526
rect 27712 40462 27764 40468
rect 27988 40520 28040 40526
rect 27988 40462 28040 40468
rect 26976 40180 27028 40186
rect 26976 40122 27028 40128
rect 28000 40050 28028 40462
rect 27988 40044 28040 40050
rect 27988 39986 28040 39992
rect 25412 38956 25464 38962
rect 25412 38898 25464 38904
rect 25780 38956 25832 38962
rect 25780 38898 25832 38904
rect 26056 38956 26108 38962
rect 26056 38898 26108 38904
rect 24860 37936 24912 37942
rect 24860 37878 24912 37884
rect 25320 37936 25372 37942
rect 25320 37878 25372 37884
rect 24124 37868 24176 37874
rect 24124 37810 24176 37816
rect 24216 37868 24268 37874
rect 24216 37810 24268 37816
rect 24136 37194 24164 37810
rect 24768 37664 24820 37670
rect 24768 37606 24820 37612
rect 24780 37330 24808 37606
rect 24768 37324 24820 37330
rect 24768 37266 24820 37272
rect 25228 37324 25280 37330
rect 25228 37266 25280 37272
rect 24124 37188 24176 37194
rect 24124 37130 24176 37136
rect 24952 36780 25004 36786
rect 24952 36722 25004 36728
rect 24676 36304 24728 36310
rect 24676 36246 24728 36252
rect 24400 36168 24452 36174
rect 24400 36110 24452 36116
rect 24308 36032 24360 36038
rect 24308 35974 24360 35980
rect 24032 35828 24084 35834
rect 24032 35770 24084 35776
rect 23848 35692 23900 35698
rect 23848 35634 23900 35640
rect 23676 35550 23796 35578
rect 23388 35158 23440 35164
rect 23570 35184 23626 35193
rect 23400 31890 23428 35158
rect 23570 35119 23626 35128
rect 23480 35012 23532 35018
rect 23480 34954 23532 34960
rect 23492 34610 23520 34954
rect 23584 34610 23612 35119
rect 23480 34604 23532 34610
rect 23480 34546 23532 34552
rect 23572 34604 23624 34610
rect 23572 34546 23624 34552
rect 23676 32910 23704 35550
rect 23756 35488 23808 35494
rect 23756 35430 23808 35436
rect 23768 35222 23796 35430
rect 23756 35216 23808 35222
rect 23756 35158 23808 35164
rect 23860 35086 23888 35634
rect 24320 35562 24348 35974
rect 24412 35698 24440 36110
rect 24584 36100 24636 36106
rect 24584 36042 24636 36048
rect 24492 35760 24544 35766
rect 24492 35702 24544 35708
rect 24400 35692 24452 35698
rect 24400 35634 24452 35640
rect 24308 35556 24360 35562
rect 24308 35498 24360 35504
rect 23848 35080 23900 35086
rect 23848 35022 23900 35028
rect 23860 34746 23888 35022
rect 23848 34740 23900 34746
rect 23848 34682 23900 34688
rect 24320 34610 24348 35498
rect 24308 34604 24360 34610
rect 24308 34546 24360 34552
rect 24504 34474 24532 35702
rect 24596 35630 24624 36042
rect 24584 35624 24636 35630
rect 24584 35566 24636 35572
rect 24596 35222 24624 35566
rect 24584 35216 24636 35222
rect 24584 35158 24636 35164
rect 24688 34610 24716 36246
rect 24860 36032 24912 36038
rect 24860 35974 24912 35980
rect 24872 35630 24900 35974
rect 24964 35698 24992 36722
rect 24952 35692 25004 35698
rect 24952 35634 25004 35640
rect 24860 35624 24912 35630
rect 24860 35566 24912 35572
rect 24768 35488 24820 35494
rect 24768 35430 24820 35436
rect 24860 35488 24912 35494
rect 24860 35430 24912 35436
rect 24780 34610 24808 35430
rect 24872 35290 24900 35430
rect 24860 35284 24912 35290
rect 24860 35226 24912 35232
rect 24872 35154 24900 35226
rect 24860 35148 24912 35154
rect 24860 35090 24912 35096
rect 24872 35034 24900 35090
rect 25044 35080 25096 35086
rect 24872 35006 24992 35034
rect 25044 35022 25096 35028
rect 24860 34944 24912 34950
rect 24860 34886 24912 34892
rect 24676 34604 24728 34610
rect 24676 34546 24728 34552
rect 24768 34604 24820 34610
rect 24768 34546 24820 34552
rect 24872 34542 24900 34886
rect 24860 34536 24912 34542
rect 24860 34478 24912 34484
rect 24492 34468 24544 34474
rect 24492 34410 24544 34416
rect 24504 33998 24532 34410
rect 24492 33992 24544 33998
rect 24492 33934 24544 33940
rect 23664 32904 23716 32910
rect 23584 32852 23664 32858
rect 23584 32846 23716 32852
rect 23584 32830 23704 32846
rect 23584 32570 23612 32830
rect 23664 32768 23716 32774
rect 23664 32710 23716 32716
rect 23572 32564 23624 32570
rect 23572 32506 23624 32512
rect 23388 31884 23440 31890
rect 23388 31826 23440 31832
rect 23676 31754 23704 32710
rect 23940 32224 23992 32230
rect 23940 32166 23992 32172
rect 23952 31822 23980 32166
rect 23940 31816 23992 31822
rect 23940 31758 23992 31764
rect 23664 31748 23716 31754
rect 23664 31690 23716 31696
rect 24504 30870 24532 33934
rect 24872 32434 24900 34478
rect 24964 33998 24992 35006
rect 25056 34610 25084 35022
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 25056 34066 25084 34546
rect 25044 34060 25096 34066
rect 25044 34002 25096 34008
rect 24952 33992 25004 33998
rect 24952 33934 25004 33940
rect 24860 32428 24912 32434
rect 24860 32370 24912 32376
rect 24584 31816 24636 31822
rect 24584 31758 24636 31764
rect 25044 31816 25096 31822
rect 25044 31758 25096 31764
rect 24492 30864 24544 30870
rect 24492 30806 24544 30812
rect 24504 30666 24532 30806
rect 24492 30660 24544 30666
rect 24492 30602 24544 30608
rect 23296 30592 23348 30598
rect 23296 30534 23348 30540
rect 24596 30258 24624 31758
rect 24768 31340 24820 31346
rect 24768 31282 24820 31288
rect 24780 30734 24808 31282
rect 24768 30728 24820 30734
rect 24768 30670 24820 30676
rect 25056 30258 25084 31758
rect 25240 31482 25268 37266
rect 25332 37262 25360 37878
rect 25424 37670 25452 38898
rect 25872 38752 25924 38758
rect 25872 38694 25924 38700
rect 25412 37664 25464 37670
rect 25412 37606 25464 37612
rect 25320 37256 25372 37262
rect 25372 37216 25452 37244
rect 25320 37198 25372 37204
rect 25320 37120 25372 37126
rect 25320 37062 25372 37068
rect 25332 36786 25360 37062
rect 25424 36854 25452 37216
rect 25688 37188 25740 37194
rect 25688 37130 25740 37136
rect 25412 36848 25464 36854
rect 25412 36790 25464 36796
rect 25320 36780 25372 36786
rect 25320 36722 25372 36728
rect 25700 35698 25728 37130
rect 25884 36174 25912 38694
rect 26068 38486 26096 38898
rect 26056 38480 26108 38486
rect 26056 38422 26108 38428
rect 28000 38350 28028 39986
rect 28356 39432 28408 39438
rect 28356 39374 28408 39380
rect 28368 39098 28396 39374
rect 28356 39092 28408 39098
rect 28356 39034 28408 39040
rect 27988 38344 28040 38350
rect 27988 38286 28040 38292
rect 27712 38276 27764 38282
rect 27712 38218 27764 38224
rect 27528 38208 27580 38214
rect 27528 38150 27580 38156
rect 27540 37942 27568 38150
rect 27724 38010 27752 38218
rect 27712 38004 27764 38010
rect 27712 37946 27764 37952
rect 27528 37936 27580 37942
rect 27528 37878 27580 37884
rect 26792 37868 26844 37874
rect 26792 37810 26844 37816
rect 27344 37868 27396 37874
rect 27344 37810 27396 37816
rect 26240 37256 26292 37262
rect 26240 37198 26292 37204
rect 26252 36854 26280 37198
rect 26240 36848 26292 36854
rect 26240 36790 26292 36796
rect 26056 36644 26108 36650
rect 26056 36586 26108 36592
rect 25872 36168 25924 36174
rect 25872 36110 25924 36116
rect 25688 35692 25740 35698
rect 25688 35634 25740 35640
rect 25884 35494 25912 36110
rect 25872 35488 25924 35494
rect 25872 35430 25924 35436
rect 25778 35184 25834 35193
rect 25778 35119 25780 35128
rect 25832 35119 25834 35128
rect 25780 35090 25832 35096
rect 25688 35080 25740 35086
rect 25688 35022 25740 35028
rect 25320 34400 25372 34406
rect 25320 34342 25372 34348
rect 25332 33522 25360 34342
rect 25700 34202 25728 35022
rect 26068 34950 26096 36586
rect 26608 36576 26660 36582
rect 26608 36518 26660 36524
rect 26240 36236 26292 36242
rect 26240 36178 26292 36184
rect 26056 34944 26108 34950
rect 26056 34886 26108 34892
rect 25688 34196 25740 34202
rect 25688 34138 25740 34144
rect 25320 33516 25372 33522
rect 25320 33458 25372 33464
rect 25412 32428 25464 32434
rect 25412 32370 25464 32376
rect 25872 32428 25924 32434
rect 25872 32370 25924 32376
rect 25424 31482 25452 32370
rect 25780 32360 25832 32366
rect 25780 32302 25832 32308
rect 25792 31482 25820 32302
rect 25228 31476 25280 31482
rect 25228 31418 25280 31424
rect 25412 31476 25464 31482
rect 25412 31418 25464 31424
rect 25780 31476 25832 31482
rect 25780 31418 25832 31424
rect 25504 31136 25556 31142
rect 25504 31078 25556 31084
rect 25516 30734 25544 31078
rect 25884 30938 25912 32370
rect 26252 32026 26280 36178
rect 26424 35216 26476 35222
rect 26424 35158 26476 35164
rect 26332 34944 26384 34950
rect 26332 34886 26384 34892
rect 26344 34678 26372 34886
rect 26332 34672 26384 34678
rect 26332 34614 26384 34620
rect 26436 34610 26464 35158
rect 26620 34610 26648 36518
rect 26424 34604 26476 34610
rect 26424 34546 26476 34552
rect 26608 34604 26660 34610
rect 26608 34546 26660 34552
rect 26424 34468 26476 34474
rect 26424 34410 26476 34416
rect 26436 33318 26464 34410
rect 26804 34066 26832 37810
rect 27252 37732 27304 37738
rect 27252 37674 27304 37680
rect 27264 37466 27292 37674
rect 27252 37460 27304 37466
rect 27252 37402 27304 37408
rect 27068 37324 27120 37330
rect 27068 37266 27120 37272
rect 26976 36848 27028 36854
rect 26976 36790 27028 36796
rect 26988 36310 27016 36790
rect 27080 36786 27108 37266
rect 27160 37256 27212 37262
rect 27160 37198 27212 37204
rect 27172 36922 27200 37198
rect 27160 36916 27212 36922
rect 27160 36858 27212 36864
rect 27068 36780 27120 36786
rect 27068 36722 27120 36728
rect 26976 36304 27028 36310
rect 26976 36246 27028 36252
rect 27080 35290 27108 36722
rect 27356 36582 27384 37810
rect 27540 37398 27568 37878
rect 27528 37392 27580 37398
rect 27528 37334 27580 37340
rect 27344 36576 27396 36582
rect 27344 36518 27396 36524
rect 27540 36174 27568 37334
rect 27712 37256 27764 37262
rect 27712 37198 27764 37204
rect 27160 36168 27212 36174
rect 27160 36110 27212 36116
rect 27528 36168 27580 36174
rect 27528 36110 27580 36116
rect 27172 35766 27200 36110
rect 27160 35760 27212 35766
rect 27160 35702 27212 35708
rect 27068 35284 27120 35290
rect 27068 35226 27120 35232
rect 27172 35154 27200 35702
rect 27724 35698 27752 37198
rect 28080 35760 28132 35766
rect 28080 35702 28132 35708
rect 27712 35692 27764 35698
rect 27712 35634 27764 35640
rect 27160 35148 27212 35154
rect 27160 35090 27212 35096
rect 27528 35080 27580 35086
rect 27528 35022 27580 35028
rect 27436 34944 27488 34950
rect 27436 34886 27488 34892
rect 26976 34740 27028 34746
rect 26976 34682 27028 34688
rect 26884 34400 26936 34406
rect 26884 34342 26936 34348
rect 26792 34060 26844 34066
rect 26792 34002 26844 34008
rect 26896 33998 26924 34342
rect 26988 33998 27016 34682
rect 27344 34604 27396 34610
rect 27344 34546 27396 34552
rect 26884 33992 26936 33998
rect 26884 33934 26936 33940
rect 26976 33992 27028 33998
rect 26976 33934 27028 33940
rect 26988 33318 27016 33934
rect 27356 33658 27384 34546
rect 27344 33652 27396 33658
rect 27344 33594 27396 33600
rect 27448 33522 27476 34886
rect 27540 33590 27568 35022
rect 27724 34610 27752 35634
rect 27896 35012 27948 35018
rect 27948 34972 28028 35000
rect 27896 34954 27948 34960
rect 27712 34604 27764 34610
rect 27712 34546 27764 34552
rect 28000 34542 28028 34972
rect 27988 34536 28040 34542
rect 27988 34478 28040 34484
rect 28092 34474 28120 35702
rect 28172 35080 28224 35086
rect 28172 35022 28224 35028
rect 28080 34468 28132 34474
rect 28080 34410 28132 34416
rect 28092 33998 28120 34410
rect 28184 34202 28212 35022
rect 28448 34604 28500 34610
rect 28448 34546 28500 34552
rect 28264 34536 28316 34542
rect 28264 34478 28316 34484
rect 28172 34196 28224 34202
rect 28172 34138 28224 34144
rect 28276 33998 28304 34478
rect 28460 33998 28488 34546
rect 28080 33992 28132 33998
rect 28080 33934 28132 33940
rect 28264 33992 28316 33998
rect 28264 33934 28316 33940
rect 28448 33992 28500 33998
rect 28448 33934 28500 33940
rect 27528 33584 27580 33590
rect 27528 33526 27580 33532
rect 27436 33516 27488 33522
rect 27436 33458 27488 33464
rect 26424 33312 26476 33318
rect 26424 33254 26476 33260
rect 26976 33312 27028 33318
rect 26976 33254 27028 33260
rect 26240 32020 26292 32026
rect 26240 31962 26292 31968
rect 26056 31680 26108 31686
rect 26056 31622 26108 31628
rect 26068 31482 26096 31622
rect 26056 31476 26108 31482
rect 26056 31418 26108 31424
rect 26056 31340 26108 31346
rect 26056 31282 26108 31288
rect 25872 30932 25924 30938
rect 25872 30874 25924 30880
rect 25504 30728 25556 30734
rect 25504 30670 25556 30676
rect 24584 30252 24636 30258
rect 24584 30194 24636 30200
rect 25044 30252 25096 30258
rect 25044 30194 25096 30200
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 24860 29504 24912 29510
rect 24860 29446 24912 29452
rect 22836 28960 22888 28966
rect 22836 28902 22888 28908
rect 22744 28756 22796 28762
rect 22744 28698 22796 28704
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22848 28558 22876 28902
rect 23308 28558 23336 29446
rect 24872 29306 24900 29446
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 23480 28620 23532 28626
rect 23480 28562 23532 28568
rect 22836 28552 22888 28558
rect 22836 28494 22888 28500
rect 23020 28552 23072 28558
rect 23020 28494 23072 28500
rect 23112 28552 23164 28558
rect 23112 28494 23164 28500
rect 23296 28552 23348 28558
rect 23296 28494 23348 28500
rect 21916 28144 21968 28150
rect 21916 28086 21968 28092
rect 21824 26988 21876 26994
rect 21928 26976 21956 28086
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22192 28008 22244 28014
rect 22192 27950 22244 27956
rect 22008 27872 22060 27878
rect 22008 27814 22060 27820
rect 22020 27538 22048 27814
rect 22204 27674 22232 27950
rect 22192 27668 22244 27674
rect 22192 27610 22244 27616
rect 22008 27532 22060 27538
rect 22008 27474 22060 27480
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 22008 26988 22060 26994
rect 21928 26948 22008 26976
rect 21824 26930 21876 26936
rect 22008 26930 22060 26936
rect 22112 26858 22140 27406
rect 22204 26976 22232 27610
rect 22296 27606 22324 28018
rect 22284 27600 22336 27606
rect 22284 27542 22336 27548
rect 22376 27056 22428 27062
rect 22376 26998 22428 27004
rect 22284 26988 22336 26994
rect 22204 26948 22284 26976
rect 22284 26930 22336 26936
rect 22100 26852 22152 26858
rect 22100 26794 22152 26800
rect 22008 26784 22060 26790
rect 22008 26726 22060 26732
rect 21824 26308 21876 26314
rect 21824 26250 21876 26256
rect 21836 25906 21864 26250
rect 22020 26246 22048 26726
rect 22008 26240 22060 26246
rect 22008 26182 22060 26188
rect 22020 25906 22048 26182
rect 21824 25900 21876 25906
rect 21824 25842 21876 25848
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 22020 25362 22048 25842
rect 22008 25356 22060 25362
rect 22008 25298 22060 25304
rect 22192 24608 22244 24614
rect 22192 24550 22244 24556
rect 22204 24342 22232 24550
rect 22192 24336 22244 24342
rect 22192 24278 22244 24284
rect 22296 24274 22324 26930
rect 22284 24268 22336 24274
rect 22284 24210 22336 24216
rect 22008 24064 22060 24070
rect 22008 24006 22060 24012
rect 22020 23866 22048 24006
rect 22008 23860 22060 23866
rect 22008 23802 22060 23808
rect 22020 23118 22048 23802
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22112 23118 22140 23666
rect 22008 23112 22060 23118
rect 22008 23054 22060 23060
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 22020 21554 22048 22918
rect 22388 22710 22416 26998
rect 22744 26308 22796 26314
rect 22744 26250 22796 26256
rect 22756 26042 22784 26250
rect 22744 26036 22796 26042
rect 22744 25978 22796 25984
rect 22848 25770 22876 28494
rect 23032 27402 23060 28494
rect 23124 28218 23152 28494
rect 23112 28212 23164 28218
rect 23112 28154 23164 28160
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 23020 27396 23072 27402
rect 23020 27338 23072 27344
rect 22928 26784 22980 26790
rect 22928 26726 22980 26732
rect 22940 25906 22968 26726
rect 23032 25906 23060 27338
rect 23216 26994 23244 27406
rect 23204 26988 23256 26994
rect 23204 26930 23256 26936
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 23400 26518 23428 26862
rect 23388 26512 23440 26518
rect 23388 26454 23440 26460
rect 22928 25900 22980 25906
rect 22928 25842 22980 25848
rect 23020 25900 23072 25906
rect 23020 25842 23072 25848
rect 23400 25838 23428 26454
rect 23492 26382 23520 28562
rect 24768 28484 24820 28490
rect 24768 28426 24820 28432
rect 24780 28218 24808 28426
rect 24768 28212 24820 28218
rect 24768 28154 24820 28160
rect 24308 28008 24360 28014
rect 24308 27950 24360 27956
rect 23480 26376 23532 26382
rect 23480 26318 23532 26324
rect 23388 25832 23440 25838
rect 23388 25774 23440 25780
rect 22836 25764 22888 25770
rect 22836 25706 22888 25712
rect 23112 25764 23164 25770
rect 23112 25706 23164 25712
rect 22652 24064 22704 24070
rect 22652 24006 22704 24012
rect 22664 23798 22692 24006
rect 22652 23792 22704 23798
rect 22652 23734 22704 23740
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 23124 22642 23152 25706
rect 23112 22636 23164 22642
rect 23112 22578 23164 22584
rect 23296 22568 23348 22574
rect 23296 22510 23348 22516
rect 22284 22432 22336 22438
rect 22284 22374 22336 22380
rect 22468 22432 22520 22438
rect 22468 22374 22520 22380
rect 22296 21622 22324 22374
rect 22480 22030 22508 22374
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22468 22024 22520 22030
rect 22468 21966 22520 21972
rect 22652 22024 22704 22030
rect 22652 21966 22704 21972
rect 22284 21616 22336 21622
rect 22284 21558 22336 21564
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 22100 21548 22152 21554
rect 22100 21490 22152 21496
rect 22112 20534 22140 21490
rect 22100 20528 22152 20534
rect 22100 20470 22152 20476
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 21836 19854 21864 20198
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 22296 19446 22324 21558
rect 22388 19922 22416 21966
rect 22480 21486 22508 21966
rect 22560 21888 22612 21894
rect 22560 21830 22612 21836
rect 22572 21554 22600 21830
rect 22664 21690 22692 21966
rect 22652 21684 22704 21690
rect 22652 21626 22704 21632
rect 22560 21548 22612 21554
rect 22560 21490 22612 21496
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22664 21010 22692 21626
rect 22928 21412 22980 21418
rect 22928 21354 22980 21360
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22836 20528 22888 20534
rect 22836 20470 22888 20476
rect 22940 20482 22968 21354
rect 23308 21010 23336 22510
rect 23400 22030 23428 25774
rect 24320 23730 24348 27950
rect 24952 26784 25004 26790
rect 24952 26726 25004 26732
rect 24964 26382 24992 26726
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 24952 26376 25004 26382
rect 24952 26318 25004 26324
rect 24412 25362 24440 26318
rect 25056 25906 25084 30194
rect 25516 29850 25544 30670
rect 26068 29850 26096 31282
rect 25504 29844 25556 29850
rect 25504 29786 25556 29792
rect 26056 29844 26108 29850
rect 26056 29786 26108 29792
rect 25504 29640 25556 29646
rect 25504 29582 25556 29588
rect 25964 29640 26016 29646
rect 25964 29582 26016 29588
rect 25412 29300 25464 29306
rect 25412 29242 25464 29248
rect 25320 29164 25372 29170
rect 25320 29106 25372 29112
rect 25136 28960 25188 28966
rect 25136 28902 25188 28908
rect 25148 28014 25176 28902
rect 25332 28150 25360 29106
rect 25320 28144 25372 28150
rect 25320 28086 25372 28092
rect 25136 28008 25188 28014
rect 25136 27950 25188 27956
rect 25332 26790 25360 28086
rect 25424 27878 25452 29242
rect 25516 29238 25544 29582
rect 25976 29306 26004 29582
rect 25964 29300 26016 29306
rect 25964 29242 26016 29248
rect 25504 29232 25556 29238
rect 25504 29174 25556 29180
rect 25516 28762 25544 29174
rect 25504 28756 25556 28762
rect 25504 28698 25556 28704
rect 25516 28150 25544 28698
rect 25504 28144 25556 28150
rect 25504 28086 25556 28092
rect 25412 27872 25464 27878
rect 25412 27814 25464 27820
rect 25424 26994 25452 27814
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 26160 26994 26188 27406
rect 26252 27062 26280 31962
rect 26332 31340 26384 31346
rect 26332 31282 26384 31288
rect 26344 30326 26372 31282
rect 26436 30666 26464 33254
rect 27528 32496 27580 32502
rect 27528 32438 27580 32444
rect 27160 32224 27212 32230
rect 27160 32166 27212 32172
rect 27172 31346 27200 32166
rect 27344 31952 27396 31958
rect 27344 31894 27396 31900
rect 27356 31822 27384 31894
rect 27344 31816 27396 31822
rect 27344 31758 27396 31764
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 27436 31136 27488 31142
rect 27436 31078 27488 31084
rect 27448 30734 27476 31078
rect 27540 30938 27568 32438
rect 28276 32298 28304 33934
rect 28460 32366 28488 33934
rect 28540 33856 28592 33862
rect 28540 33798 28592 33804
rect 28448 32360 28500 32366
rect 28448 32302 28500 32308
rect 27896 32292 27948 32298
rect 27896 32234 27948 32240
rect 28264 32292 28316 32298
rect 28264 32234 28316 32240
rect 27528 30932 27580 30938
rect 27528 30874 27580 30880
rect 26976 30728 27028 30734
rect 26976 30670 27028 30676
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 26424 30660 26476 30666
rect 26424 30602 26476 30608
rect 26608 30592 26660 30598
rect 26608 30534 26660 30540
rect 26332 30320 26384 30326
rect 26332 30262 26384 30268
rect 26240 27056 26292 27062
rect 26240 26998 26292 27004
rect 25412 26988 25464 26994
rect 25412 26930 25464 26936
rect 25872 26988 25924 26994
rect 25872 26930 25924 26936
rect 26148 26988 26200 26994
rect 26148 26930 26200 26936
rect 25884 26790 25912 26930
rect 26056 26920 26108 26926
rect 26056 26862 26108 26868
rect 25320 26784 25372 26790
rect 25320 26726 25372 26732
rect 25872 26784 25924 26790
rect 25872 26726 25924 26732
rect 25044 25900 25096 25906
rect 25044 25842 25096 25848
rect 25056 25498 25084 25842
rect 25332 25838 25360 26726
rect 26068 26586 26096 26862
rect 26056 26580 26108 26586
rect 26056 26522 26108 26528
rect 26620 26364 26648 30534
rect 26988 29850 27016 30670
rect 27540 30394 27568 30874
rect 27528 30388 27580 30394
rect 27528 30330 27580 30336
rect 27908 30122 27936 32234
rect 28356 32224 28408 32230
rect 28356 32166 28408 32172
rect 28080 31340 28132 31346
rect 28080 31282 28132 31288
rect 28092 30734 28120 31282
rect 28368 30734 28396 32166
rect 28552 31414 28580 33798
rect 28632 32292 28684 32298
rect 28632 32234 28684 32240
rect 28540 31408 28592 31414
rect 28540 31350 28592 31356
rect 28644 30870 28672 32234
rect 28632 30864 28684 30870
rect 28632 30806 28684 30812
rect 28080 30728 28132 30734
rect 28080 30670 28132 30676
rect 28356 30728 28408 30734
rect 28356 30670 28408 30676
rect 28264 30252 28316 30258
rect 28264 30194 28316 30200
rect 27896 30116 27948 30122
rect 27896 30058 27948 30064
rect 26976 29844 27028 29850
rect 26976 29786 27028 29792
rect 27160 29708 27212 29714
rect 27160 29650 27212 29656
rect 26884 29640 26936 29646
rect 26884 29582 26936 29588
rect 26896 29306 26924 29582
rect 26884 29300 26936 29306
rect 26884 29242 26936 29248
rect 26896 28558 26924 29242
rect 26884 28552 26936 28558
rect 26884 28494 26936 28500
rect 27068 28552 27120 28558
rect 27068 28494 27120 28500
rect 26896 28082 26924 28494
rect 27080 28082 27108 28494
rect 26884 28076 26936 28082
rect 26884 28018 26936 28024
rect 27068 28076 27120 28082
rect 27068 28018 27120 28024
rect 27172 28014 27200 29650
rect 27620 29164 27672 29170
rect 27620 29106 27672 29112
rect 27632 28762 27660 29106
rect 27620 28756 27672 28762
rect 27620 28698 27672 28704
rect 27252 28552 27304 28558
rect 27252 28494 27304 28500
rect 27264 28218 27292 28494
rect 27252 28212 27304 28218
rect 27252 28154 27304 28160
rect 27160 28008 27212 28014
rect 27160 27950 27212 27956
rect 27344 27600 27396 27606
rect 27344 27542 27396 27548
rect 27356 26994 27384 27542
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27724 26994 27752 27406
rect 27804 27396 27856 27402
rect 27804 27338 27856 27344
rect 27344 26988 27396 26994
rect 27344 26930 27396 26936
rect 27712 26988 27764 26994
rect 27712 26930 27764 26936
rect 27620 26920 27672 26926
rect 27816 26874 27844 27338
rect 27672 26868 27844 26874
rect 27620 26862 27844 26868
rect 26700 26852 26752 26858
rect 27632 26846 27844 26862
rect 26700 26794 26752 26800
rect 26712 26518 26740 26794
rect 27160 26784 27212 26790
rect 27160 26726 27212 26732
rect 26700 26512 26752 26518
rect 26700 26454 26752 26460
rect 26620 26336 26740 26364
rect 25320 25832 25372 25838
rect 25320 25774 25372 25780
rect 25044 25492 25096 25498
rect 25044 25434 25096 25440
rect 24400 25356 24452 25362
rect 24400 25298 24452 25304
rect 24492 25220 24544 25226
rect 24492 25162 24544 25168
rect 24504 24954 24532 25162
rect 24492 24948 24544 24954
rect 24492 24890 24544 24896
rect 25332 24818 25360 25774
rect 25320 24812 25372 24818
rect 25320 24754 25372 24760
rect 25688 24744 25740 24750
rect 25688 24686 25740 24692
rect 25700 24274 25728 24686
rect 25688 24268 25740 24274
rect 25688 24210 25740 24216
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 25044 23656 25096 23662
rect 25044 23598 25096 23604
rect 25056 23118 25084 23598
rect 25044 23112 25096 23118
rect 25044 23054 25096 23060
rect 24676 23044 24728 23050
rect 24676 22986 24728 22992
rect 24688 22778 24716 22986
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24952 22704 25004 22710
rect 24952 22646 25004 22652
rect 24216 22432 24268 22438
rect 24216 22374 24268 22380
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 24228 21554 24256 22374
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 23296 21004 23348 21010
rect 23296 20946 23348 20952
rect 23308 20534 23336 20946
rect 23296 20528 23348 20534
rect 22848 19922 22876 20470
rect 22940 20466 23060 20482
rect 23296 20470 23348 20476
rect 22940 20460 23072 20466
rect 22940 20454 23020 20460
rect 22940 20262 22968 20454
rect 23020 20402 23072 20408
rect 23020 20324 23072 20330
rect 23020 20266 23072 20272
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 22376 19916 22428 19922
rect 22376 19858 22428 19864
rect 22836 19916 22888 19922
rect 22836 19858 22888 19864
rect 22388 19514 22416 19858
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22284 19440 22336 19446
rect 22284 19382 22336 19388
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22112 18970 22140 19314
rect 22848 18970 22876 19858
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 22836 18964 22888 18970
rect 22836 18906 22888 18912
rect 22848 18766 22876 18906
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 23032 18698 23060 20266
rect 23020 18692 23072 18698
rect 23020 18634 23072 18640
rect 23308 18630 23336 20470
rect 23388 20460 23440 20466
rect 23388 20402 23440 20408
rect 23400 19514 23428 20402
rect 23572 20256 23624 20262
rect 23572 20198 23624 20204
rect 23584 19990 23612 20198
rect 23572 19984 23624 19990
rect 23572 19926 23624 19932
rect 24964 19854 24992 22646
rect 25056 21554 25084 23054
rect 25700 22710 25728 24210
rect 26608 24132 26660 24138
rect 26608 24074 26660 24080
rect 25964 24064 26016 24070
rect 25964 24006 26016 24012
rect 25976 23798 26004 24006
rect 25964 23792 26016 23798
rect 25964 23734 26016 23740
rect 26620 23662 26648 24074
rect 26608 23656 26660 23662
rect 26608 23598 26660 23604
rect 25780 22976 25832 22982
rect 25780 22918 25832 22924
rect 25688 22704 25740 22710
rect 25688 22646 25740 22652
rect 25792 22642 25820 22918
rect 25780 22636 25832 22642
rect 25780 22578 25832 22584
rect 26712 22098 26740 26336
rect 27172 26314 27200 26726
rect 27816 26586 27844 26846
rect 27804 26580 27856 26586
rect 27804 26522 27856 26528
rect 27160 26308 27212 26314
rect 27160 26250 27212 26256
rect 27344 24812 27396 24818
rect 27344 24754 27396 24760
rect 27356 24342 27384 24754
rect 27344 24336 27396 24342
rect 27344 24278 27396 24284
rect 26792 24200 26844 24206
rect 26792 24142 26844 24148
rect 26976 24200 27028 24206
rect 26976 24142 27028 24148
rect 26804 23322 26832 24142
rect 26988 23730 27016 24142
rect 27356 24070 27384 24278
rect 27344 24064 27396 24070
rect 27344 24006 27396 24012
rect 27356 23866 27384 24006
rect 27344 23860 27396 23866
rect 27344 23802 27396 23808
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 26792 23316 26844 23322
rect 26792 23258 26844 23264
rect 26804 22234 26832 23258
rect 26988 22982 27016 23666
rect 27356 23322 27384 23802
rect 27908 23730 27936 30058
rect 28276 28762 28304 30194
rect 28736 29238 28764 45902
rect 29288 45558 29316 46922
rect 29564 46170 29592 46990
rect 30932 46368 30984 46374
rect 30932 46310 30984 46316
rect 29552 46164 29604 46170
rect 29552 46106 29604 46112
rect 30944 46034 30972 46310
rect 31588 46034 31616 49200
rect 32232 47138 32260 49200
rect 35806 49056 35862 49065
rect 35806 48991 35862 49000
rect 35346 47696 35402 47705
rect 35346 47631 35402 47640
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 32232 47122 32352 47138
rect 32232 47116 32364 47122
rect 32232 47110 32312 47116
rect 32312 47058 32364 47064
rect 32128 47048 32180 47054
rect 32128 46990 32180 46996
rect 32140 46578 32168 46990
rect 32312 46980 32364 46986
rect 32312 46922 32364 46928
rect 32128 46572 32180 46578
rect 32128 46514 32180 46520
rect 30932 46028 30984 46034
rect 30932 45970 30984 45976
rect 31576 46028 31628 46034
rect 31576 45970 31628 45976
rect 31116 45892 31168 45898
rect 31116 45834 31168 45840
rect 31128 45626 31156 45834
rect 31116 45620 31168 45626
rect 31116 45562 31168 45568
rect 32324 45558 32352 46922
rect 35360 46646 35388 47631
rect 33232 46640 33284 46646
rect 33232 46582 33284 46588
rect 35348 46640 35400 46646
rect 35348 46582 35400 46588
rect 33244 45966 33272 46582
rect 35820 46510 35848 48991
rect 35912 47462 35940 49422
rect 36054 49200 36166 49422
rect 37342 49200 37454 50000
rect 37986 49314 38098 50000
rect 37986 49286 38240 49314
rect 37986 49200 38098 49286
rect 35900 47456 35952 47462
rect 35900 47398 35952 47404
rect 37188 47456 37240 47462
rect 37188 47398 37240 47404
rect 36728 47116 36780 47122
rect 36728 47058 36780 47064
rect 36452 47048 36504 47054
rect 36452 46990 36504 46996
rect 33324 46504 33376 46510
rect 33324 46446 33376 46452
rect 35808 46504 35860 46510
rect 35808 46446 35860 46452
rect 33336 46170 33364 46446
rect 33876 46436 33928 46442
rect 33876 46378 33928 46384
rect 33888 46170 33916 46378
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 33324 46164 33376 46170
rect 33324 46106 33376 46112
rect 33876 46164 33928 46170
rect 33876 46106 33928 46112
rect 36464 46034 36492 46990
rect 36740 46578 36768 47058
rect 36728 46572 36780 46578
rect 36728 46514 36780 46520
rect 37094 46336 37150 46345
rect 37094 46271 37150 46280
rect 36452 46028 36504 46034
rect 36452 45970 36504 45976
rect 33232 45960 33284 45966
rect 33232 45902 33284 45908
rect 35806 45656 35862 45665
rect 35806 45591 35862 45600
rect 29276 45552 29328 45558
rect 29276 45494 29328 45500
rect 32312 45552 32364 45558
rect 32312 45494 32364 45500
rect 31208 45484 31260 45490
rect 31208 45426 31260 45432
rect 32404 45484 32456 45490
rect 32404 45426 32456 45432
rect 29276 45416 29328 45422
rect 29276 45358 29328 45364
rect 29288 44266 29316 45358
rect 29920 44396 29972 44402
rect 29920 44338 29972 44344
rect 29276 44260 29328 44266
rect 29276 44202 29328 44208
rect 29288 42242 29316 44202
rect 29828 44192 29880 44198
rect 29828 44134 29880 44140
rect 29840 43790 29868 44134
rect 29828 43784 29880 43790
rect 29828 43726 29880 43732
rect 29552 43648 29604 43654
rect 29552 43590 29604 43596
rect 29564 43314 29592 43590
rect 29932 43450 29960 44338
rect 30932 43648 30984 43654
rect 30932 43590 30984 43596
rect 29920 43444 29972 43450
rect 29920 43386 29972 43392
rect 29552 43308 29604 43314
rect 30288 43308 30340 43314
rect 29604 43268 29684 43296
rect 29552 43250 29604 43256
rect 29368 42628 29420 42634
rect 29368 42570 29420 42576
rect 29380 42362 29408 42570
rect 29656 42566 29684 43268
rect 30288 43250 30340 43256
rect 29920 42696 29972 42702
rect 29920 42638 29972 42644
rect 29644 42560 29696 42566
rect 29644 42502 29696 42508
rect 29368 42356 29420 42362
rect 29368 42298 29420 42304
rect 29288 42214 29408 42242
rect 28908 41472 28960 41478
rect 28908 41414 28960 41420
rect 28920 41206 28948 41414
rect 28908 41200 28960 41206
rect 28908 41142 28960 41148
rect 28908 40044 28960 40050
rect 28908 39986 28960 39992
rect 28920 39642 28948 39986
rect 28908 39636 28960 39642
rect 28908 39578 28960 39584
rect 28908 37868 28960 37874
rect 28908 37810 28960 37816
rect 28920 36922 28948 37810
rect 29000 37800 29052 37806
rect 29000 37742 29052 37748
rect 29012 37466 29040 37742
rect 29000 37460 29052 37466
rect 29000 37402 29052 37408
rect 28908 36916 28960 36922
rect 28908 36858 28960 36864
rect 29276 36168 29328 36174
rect 29276 36110 29328 36116
rect 29092 34536 29144 34542
rect 29092 34478 29144 34484
rect 29104 34066 29132 34478
rect 29092 34060 29144 34066
rect 29092 34002 29144 34008
rect 28908 32428 28960 32434
rect 28908 32370 28960 32376
rect 28920 31822 28948 32370
rect 28908 31816 28960 31822
rect 28908 31758 28960 31764
rect 28920 30326 28948 31758
rect 29288 31482 29316 36110
rect 29276 31476 29328 31482
rect 29276 31418 29328 31424
rect 28908 30320 28960 30326
rect 28908 30262 28960 30268
rect 28816 30252 28868 30258
rect 28816 30194 28868 30200
rect 29000 30252 29052 30258
rect 29000 30194 29052 30200
rect 28724 29232 28776 29238
rect 28724 29174 28776 29180
rect 28264 28756 28316 28762
rect 28264 28698 28316 28704
rect 28172 28484 28224 28490
rect 28172 28426 28224 28432
rect 28184 28082 28212 28426
rect 28276 28218 28304 28698
rect 28828 28490 28856 30194
rect 29012 29850 29040 30194
rect 29000 29844 29052 29850
rect 29000 29786 29052 29792
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 29276 29640 29328 29646
rect 29276 29582 29328 29588
rect 28920 29238 28948 29582
rect 28908 29232 28960 29238
rect 28908 29174 28960 29180
rect 28920 28762 28948 29174
rect 29288 29102 29316 29582
rect 29380 29578 29408 42214
rect 29656 42022 29684 42502
rect 29932 42294 29960 42638
rect 30012 42628 30064 42634
rect 30012 42570 30064 42576
rect 29920 42288 29972 42294
rect 29920 42230 29972 42236
rect 29644 42016 29696 42022
rect 29644 41958 29696 41964
rect 29932 41682 29960 42230
rect 30024 42158 30052 42570
rect 30012 42152 30064 42158
rect 30012 42094 30064 42100
rect 30300 42106 30328 43250
rect 30944 42770 30972 43590
rect 31116 43308 31168 43314
rect 31116 43250 31168 43256
rect 30380 42764 30432 42770
rect 30380 42706 30432 42712
rect 30932 42764 30984 42770
rect 30932 42706 30984 42712
rect 30392 42226 30420 42706
rect 31128 42362 31156 43250
rect 31116 42356 31168 42362
rect 31116 42298 31168 42304
rect 30380 42220 30432 42226
rect 30380 42162 30432 42168
rect 30472 42220 30524 42226
rect 30472 42162 30524 42168
rect 30484 42106 30512 42162
rect 29920 41676 29972 41682
rect 29920 41618 29972 41624
rect 30024 41274 30052 42094
rect 30300 42078 30512 42106
rect 30392 41614 30420 42078
rect 31220 41682 31248 45426
rect 31944 43104 31996 43110
rect 31944 43046 31996 43052
rect 31956 42702 31984 43046
rect 31944 42696 31996 42702
rect 31944 42638 31996 42644
rect 31208 41676 31260 41682
rect 31208 41618 31260 41624
rect 30380 41608 30432 41614
rect 30380 41550 30432 41556
rect 31116 41608 31168 41614
rect 31116 41550 31168 41556
rect 30012 41268 30064 41274
rect 30012 41210 30064 41216
rect 29552 39364 29604 39370
rect 29552 39306 29604 39312
rect 29564 36718 29592 39306
rect 29828 38004 29880 38010
rect 29828 37946 29880 37952
rect 29552 36712 29604 36718
rect 29552 36654 29604 36660
rect 29644 36644 29696 36650
rect 29644 36586 29696 36592
rect 29656 35154 29684 36586
rect 29552 35148 29604 35154
rect 29552 35090 29604 35096
rect 29644 35148 29696 35154
rect 29644 35090 29696 35096
rect 29564 34542 29592 35090
rect 29552 34536 29604 34542
rect 29552 34478 29604 34484
rect 29564 33998 29592 34478
rect 29552 33992 29604 33998
rect 29552 33934 29604 33940
rect 29656 33590 29684 35090
rect 29840 33862 29868 37946
rect 30104 37868 30156 37874
rect 30104 37810 30156 37816
rect 30012 37664 30064 37670
rect 30012 37606 30064 37612
rect 30024 37194 30052 37606
rect 30012 37188 30064 37194
rect 30012 37130 30064 37136
rect 30116 36922 30144 37810
rect 30104 36916 30156 36922
rect 30104 36858 30156 36864
rect 30196 36712 30248 36718
rect 30196 36654 30248 36660
rect 30208 36582 30236 36654
rect 30196 36576 30248 36582
rect 30196 36518 30248 36524
rect 30208 35154 30236 36518
rect 30196 35148 30248 35154
rect 30196 35090 30248 35096
rect 29920 35080 29972 35086
rect 29920 35022 29972 35028
rect 29932 34746 29960 35022
rect 29920 34740 29972 34746
rect 29920 34682 29972 34688
rect 29828 33856 29880 33862
rect 29828 33798 29880 33804
rect 29644 33584 29696 33590
rect 29644 33526 29696 33532
rect 29840 33318 29868 33798
rect 30392 33522 30420 41550
rect 31128 41274 31156 41550
rect 31116 41268 31168 41274
rect 31116 41210 31168 41216
rect 30932 41132 30984 41138
rect 30932 41074 30984 41080
rect 30656 40180 30708 40186
rect 30656 40122 30708 40128
rect 30668 39506 30696 40122
rect 30748 40112 30800 40118
rect 30748 40054 30800 40060
rect 30656 39500 30708 39506
rect 30656 39442 30708 39448
rect 30668 38350 30696 39442
rect 30656 38344 30708 38350
rect 30656 38286 30708 38292
rect 30760 36854 30788 40054
rect 30840 37120 30892 37126
rect 30840 37062 30892 37068
rect 30748 36848 30800 36854
rect 30748 36790 30800 36796
rect 30656 35556 30708 35562
rect 30656 35498 30708 35504
rect 30472 34944 30524 34950
rect 30472 34886 30524 34892
rect 30484 33998 30512 34886
rect 30564 34604 30616 34610
rect 30564 34546 30616 34552
rect 30576 34202 30604 34546
rect 30564 34196 30616 34202
rect 30564 34138 30616 34144
rect 30668 34134 30696 35498
rect 30656 34128 30708 34134
rect 30656 34070 30708 34076
rect 30472 33992 30524 33998
rect 30472 33934 30524 33940
rect 30668 33658 30696 34070
rect 30656 33652 30708 33658
rect 30656 33594 30708 33600
rect 30380 33516 30432 33522
rect 30380 33458 30432 33464
rect 29828 33312 29880 33318
rect 29828 33254 29880 33260
rect 30392 32910 30420 33458
rect 30380 32904 30432 32910
rect 30380 32846 30432 32852
rect 30392 32502 30420 32846
rect 30380 32496 30432 32502
rect 30380 32438 30432 32444
rect 30472 32496 30524 32502
rect 30472 32438 30524 32444
rect 29828 32360 29880 32366
rect 29828 32302 29880 32308
rect 29552 31816 29604 31822
rect 29840 31800 29868 32302
rect 30380 32224 30432 32230
rect 30380 32166 30432 32172
rect 30392 31890 30420 32166
rect 30380 31884 30432 31890
rect 30380 31826 30432 31832
rect 29920 31816 29972 31822
rect 29552 31758 29604 31764
rect 29828 31794 29880 31800
rect 29460 31680 29512 31686
rect 29460 31622 29512 31628
rect 29472 31346 29500 31622
rect 29460 31340 29512 31346
rect 29460 31282 29512 31288
rect 29564 30954 29592 31758
rect 29920 31758 29972 31764
rect 30196 31816 30248 31822
rect 30196 31758 30248 31764
rect 29828 31736 29880 31742
rect 29736 31340 29788 31346
rect 29932 31328 29960 31758
rect 30208 31498 30236 31758
rect 30484 31754 30512 32438
rect 30760 32026 30788 36790
rect 30852 36786 30880 37062
rect 30840 36780 30892 36786
rect 30840 36722 30892 36728
rect 30748 32020 30800 32026
rect 30852 32008 30880 36722
rect 30944 32570 30972 41074
rect 30932 32564 30984 32570
rect 30932 32506 30984 32512
rect 30932 32020 30984 32026
rect 30852 31980 30932 32008
rect 30748 31962 30800 31968
rect 30932 31962 30984 31968
rect 30024 31482 30236 31498
rect 30392 31726 30512 31754
rect 30392 31482 30420 31726
rect 30012 31476 30236 31482
rect 30064 31470 30236 31476
rect 30380 31476 30432 31482
rect 30012 31418 30064 31424
rect 30380 31418 30432 31424
rect 29788 31300 29960 31328
rect 29736 31282 29788 31288
rect 29472 30938 29592 30954
rect 29748 30938 29776 31282
rect 29460 30932 29592 30938
rect 29512 30926 29592 30932
rect 29736 30932 29788 30938
rect 29460 30874 29512 30880
rect 29736 30874 29788 30880
rect 30564 30320 30616 30326
rect 30564 30262 30616 30268
rect 29644 30252 29696 30258
rect 29644 30194 29696 30200
rect 29460 30048 29512 30054
rect 29460 29990 29512 29996
rect 29472 29578 29500 29990
rect 29368 29572 29420 29578
rect 29368 29514 29420 29520
rect 29460 29572 29512 29578
rect 29460 29514 29512 29520
rect 29656 29306 29684 30194
rect 30380 30048 30432 30054
rect 30380 29990 30432 29996
rect 30392 29646 30420 29990
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 29644 29300 29696 29306
rect 29644 29242 29696 29248
rect 29276 29096 29328 29102
rect 29276 29038 29328 29044
rect 30392 29034 30420 29582
rect 30576 29306 30604 30262
rect 30656 29776 30708 29782
rect 30656 29718 30708 29724
rect 30564 29300 30616 29306
rect 30564 29242 30616 29248
rect 30668 29170 30696 29718
rect 30656 29164 30708 29170
rect 30656 29106 30708 29112
rect 30380 29028 30432 29034
rect 30380 28970 30432 28976
rect 30656 29028 30708 29034
rect 30656 28970 30708 28976
rect 28908 28756 28960 28762
rect 28908 28698 28960 28704
rect 28448 28484 28500 28490
rect 28448 28426 28500 28432
rect 28816 28484 28868 28490
rect 28816 28426 28868 28432
rect 28264 28212 28316 28218
rect 28264 28154 28316 28160
rect 28172 28076 28224 28082
rect 28172 28018 28224 28024
rect 28184 27470 28212 28018
rect 28172 27464 28224 27470
rect 28172 27406 28224 27412
rect 28276 27402 28304 28154
rect 28460 28150 28488 28426
rect 28448 28144 28500 28150
rect 28448 28086 28500 28092
rect 28264 27396 28316 27402
rect 28264 27338 28316 27344
rect 28460 26858 28488 28086
rect 28920 28082 28948 28698
rect 28908 28076 28960 28082
rect 28908 28018 28960 28024
rect 30380 28076 30432 28082
rect 30380 28018 30432 28024
rect 29092 27872 29144 27878
rect 29092 27814 29144 27820
rect 29104 27062 29132 27814
rect 29092 27056 29144 27062
rect 29092 26998 29144 27004
rect 30392 26994 30420 28018
rect 30668 27334 30696 28970
rect 30760 27470 30788 31962
rect 30944 31482 30972 31962
rect 30932 31476 30984 31482
rect 30932 31418 30984 31424
rect 30932 30728 30984 30734
rect 30932 30670 30984 30676
rect 30944 29850 30972 30670
rect 30932 29844 30984 29850
rect 30932 29786 30984 29792
rect 30840 29572 30892 29578
rect 30840 29514 30892 29520
rect 30852 27606 30880 29514
rect 31220 29510 31248 41618
rect 31760 41064 31812 41070
rect 31760 41006 31812 41012
rect 31772 40050 31800 41006
rect 31576 40044 31628 40050
rect 31576 39986 31628 39992
rect 31760 40044 31812 40050
rect 31760 39986 31812 39992
rect 31392 39840 31444 39846
rect 31392 39782 31444 39788
rect 31404 38962 31432 39782
rect 31588 39642 31616 39986
rect 31576 39636 31628 39642
rect 31576 39578 31628 39584
rect 31772 39030 31800 39986
rect 32128 39840 32180 39846
rect 32128 39782 32180 39788
rect 32140 39438 32168 39782
rect 32128 39432 32180 39438
rect 32128 39374 32180 39380
rect 32312 39432 32364 39438
rect 32312 39374 32364 39380
rect 31760 39024 31812 39030
rect 31760 38966 31812 38972
rect 32140 38978 32168 39374
rect 31392 38956 31444 38962
rect 31392 38898 31444 38904
rect 31852 38956 31904 38962
rect 32140 38950 32260 38978
rect 32324 38962 32352 39374
rect 31852 38898 31904 38904
rect 31668 38344 31720 38350
rect 31668 38286 31720 38292
rect 31680 37806 31708 38286
rect 31668 37800 31720 37806
rect 31668 37742 31720 37748
rect 31864 37262 31892 38898
rect 32128 38888 32180 38894
rect 32128 38830 32180 38836
rect 32140 38418 32168 38830
rect 32128 38412 32180 38418
rect 32128 38354 32180 38360
rect 32140 37942 32168 38354
rect 32232 38282 32260 38950
rect 32312 38956 32364 38962
rect 32312 38898 32364 38904
rect 32312 38752 32364 38758
rect 32312 38694 32364 38700
rect 32324 38554 32352 38694
rect 32312 38548 32364 38554
rect 32312 38490 32364 38496
rect 32220 38276 32272 38282
rect 32220 38218 32272 38224
rect 32128 37936 32180 37942
rect 32128 37878 32180 37884
rect 31760 37256 31812 37262
rect 31760 37198 31812 37204
rect 31852 37256 31904 37262
rect 31852 37198 31904 37204
rect 31392 37120 31444 37126
rect 31392 37062 31444 37068
rect 31404 36174 31432 37062
rect 31772 36854 31800 37198
rect 31760 36848 31812 36854
rect 31760 36790 31812 36796
rect 31576 36780 31628 36786
rect 31576 36722 31628 36728
rect 31588 36310 31616 36722
rect 31576 36304 31628 36310
rect 31576 36246 31628 36252
rect 31392 36168 31444 36174
rect 31392 36110 31444 36116
rect 31864 35018 31892 37198
rect 32140 36922 32168 37878
rect 32232 37874 32260 38218
rect 32324 38010 32352 38490
rect 32312 38004 32364 38010
rect 32312 37946 32364 37952
rect 32220 37868 32272 37874
rect 32220 37810 32272 37816
rect 32324 37330 32352 37946
rect 32312 37324 32364 37330
rect 32312 37266 32364 37272
rect 32128 36916 32180 36922
rect 32128 36858 32180 36864
rect 32036 35080 32088 35086
rect 32036 35022 32088 35028
rect 31852 35012 31904 35018
rect 31852 34954 31904 34960
rect 31944 34944 31996 34950
rect 31944 34886 31996 34892
rect 31956 33862 31984 34886
rect 32048 34542 32076 35022
rect 32128 35012 32180 35018
rect 32128 34954 32180 34960
rect 32036 34536 32088 34542
rect 32036 34478 32088 34484
rect 31944 33856 31996 33862
rect 31944 33798 31996 33804
rect 31300 33448 31352 33454
rect 31300 33390 31352 33396
rect 31312 32502 31340 33390
rect 31300 32496 31352 32502
rect 31300 32438 31352 32444
rect 32048 32366 32076 34478
rect 32140 34066 32168 34954
rect 32416 34490 32444 45426
rect 35820 45422 35848 45591
rect 35808 45416 35860 45422
rect 35808 45358 35860 45364
rect 36544 45416 36596 45422
rect 36544 45358 36596 45364
rect 36728 45416 36780 45422
rect 36728 45358 36780 45364
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 36556 44538 36584 45358
rect 36544 44532 36596 44538
rect 36544 44474 36596 44480
rect 36740 44402 36768 45358
rect 37108 44946 37136 46271
rect 37096 44940 37148 44946
rect 37096 44882 37148 44888
rect 36728 44396 36780 44402
rect 36728 44338 36780 44344
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 36268 43784 36320 43790
rect 36268 43726 36320 43732
rect 36280 43314 36308 43726
rect 35808 43308 35860 43314
rect 35808 43250 35860 43256
rect 36268 43308 36320 43314
rect 36268 43250 36320 43256
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 35820 42945 35848 43250
rect 35900 43104 35952 43110
rect 35900 43046 35952 43052
rect 35806 42936 35862 42945
rect 35806 42871 35862 42880
rect 33048 42696 33100 42702
rect 33048 42638 33100 42644
rect 33060 42158 33088 42638
rect 33876 42220 33928 42226
rect 33876 42162 33928 42168
rect 33048 42152 33100 42158
rect 33048 42094 33100 42100
rect 33060 41206 33088 42094
rect 33888 41818 33916 42162
rect 34796 42016 34848 42022
rect 34796 41958 34848 41964
rect 33876 41812 33928 41818
rect 33876 41754 33928 41760
rect 34244 41608 34296 41614
rect 34244 41550 34296 41556
rect 34520 41608 34572 41614
rect 34520 41550 34572 41556
rect 34610 41576 34666 41585
rect 34256 41274 34284 41550
rect 34244 41268 34296 41274
rect 34244 41210 34296 41216
rect 33048 41200 33100 41206
rect 33048 41142 33100 41148
rect 32680 41132 32732 41138
rect 32680 41074 32732 41080
rect 32692 40730 32720 41074
rect 34532 40730 34560 41550
rect 34610 41511 34612 41520
rect 34664 41511 34666 41520
rect 34612 41482 34664 41488
rect 34808 41414 34836 41958
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34716 41386 34836 41414
rect 34716 40730 34744 41386
rect 34796 41064 34848 41070
rect 34796 41006 34848 41012
rect 35348 41064 35400 41070
rect 35348 41006 35400 41012
rect 32680 40724 32732 40730
rect 32680 40666 32732 40672
rect 34520 40724 34572 40730
rect 34520 40666 34572 40672
rect 34704 40724 34756 40730
rect 34704 40666 34756 40672
rect 34612 40588 34664 40594
rect 34612 40530 34664 40536
rect 32864 40520 32916 40526
rect 32864 40462 32916 40468
rect 32876 39642 32904 40462
rect 33600 40384 33652 40390
rect 33600 40326 33652 40332
rect 33232 40044 33284 40050
rect 33232 39986 33284 39992
rect 33244 39642 33272 39986
rect 32864 39636 32916 39642
rect 32864 39578 32916 39584
rect 33232 39636 33284 39642
rect 33232 39578 33284 39584
rect 32496 39432 32548 39438
rect 32496 39374 32548 39380
rect 32508 39098 32536 39374
rect 32496 39092 32548 39098
rect 32496 39034 32548 39040
rect 33612 38350 33640 40326
rect 34244 40044 34296 40050
rect 34244 39986 34296 39992
rect 33968 39976 34020 39982
rect 33968 39918 34020 39924
rect 33980 38962 34008 39918
rect 34256 39642 34284 39986
rect 34244 39636 34296 39642
rect 34244 39578 34296 39584
rect 34624 39370 34652 40530
rect 34716 40050 34744 40666
rect 34808 40526 34836 41006
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34796 40520 34848 40526
rect 34796 40462 34848 40468
rect 34704 40044 34756 40050
rect 34704 39986 34756 39992
rect 34716 39506 34744 39986
rect 34808 39574 34836 40462
rect 35360 40458 35388 41006
rect 35808 40928 35860 40934
rect 35808 40870 35860 40876
rect 35820 40526 35848 40870
rect 35808 40520 35860 40526
rect 35808 40462 35860 40468
rect 35348 40452 35400 40458
rect 35348 40394 35400 40400
rect 35360 39846 35388 40394
rect 35624 40384 35676 40390
rect 35624 40326 35676 40332
rect 35348 39840 35400 39846
rect 35348 39782 35400 39788
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34796 39568 34848 39574
rect 34796 39510 34848 39516
rect 34704 39500 34756 39506
rect 34704 39442 34756 39448
rect 34612 39364 34664 39370
rect 34612 39306 34664 39312
rect 35360 39302 35388 39782
rect 34704 39296 34756 39302
rect 34704 39238 34756 39244
rect 34980 39296 35032 39302
rect 34980 39238 35032 39244
rect 35348 39296 35400 39302
rect 35348 39238 35400 39244
rect 33968 38956 34020 38962
rect 33968 38898 34020 38904
rect 33600 38344 33652 38350
rect 33600 38286 33652 38292
rect 33140 38208 33192 38214
rect 33140 38150 33192 38156
rect 32772 37664 32824 37670
rect 32772 37606 32824 37612
rect 32784 37262 32812 37606
rect 33152 37262 33180 38150
rect 34520 37868 34572 37874
rect 34520 37810 34572 37816
rect 34336 37664 34388 37670
rect 34336 37606 34388 37612
rect 33232 37324 33284 37330
rect 33232 37266 33284 37272
rect 32772 37256 32824 37262
rect 32772 37198 32824 37204
rect 33140 37256 33192 37262
rect 33140 37198 33192 37204
rect 32956 37188 33008 37194
rect 32956 37130 33008 37136
rect 32588 37120 32640 37126
rect 32588 37062 32640 37068
rect 32600 34678 32628 37062
rect 32772 36916 32824 36922
rect 32772 36858 32824 36864
rect 32784 36582 32812 36858
rect 32864 36848 32916 36854
rect 32864 36790 32916 36796
rect 32876 36582 32904 36790
rect 32772 36576 32824 36582
rect 32772 36518 32824 36524
rect 32864 36576 32916 36582
rect 32864 36518 32916 36524
rect 32876 35086 32904 36518
rect 32864 35080 32916 35086
rect 32864 35022 32916 35028
rect 32588 34672 32640 34678
rect 32588 34614 32640 34620
rect 32416 34462 32628 34490
rect 32128 34060 32180 34066
rect 32128 34002 32180 34008
rect 32220 33992 32272 33998
rect 32220 33934 32272 33940
rect 32232 32910 32260 33934
rect 32404 33108 32456 33114
rect 32404 33050 32456 33056
rect 32220 32904 32272 32910
rect 32220 32846 32272 32852
rect 32232 32502 32260 32846
rect 32220 32496 32272 32502
rect 32220 32438 32272 32444
rect 32036 32360 32088 32366
rect 32036 32302 32088 32308
rect 31300 31816 31352 31822
rect 31300 31758 31352 31764
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 31312 31346 31340 31758
rect 31300 31340 31352 31346
rect 31300 31282 31352 31288
rect 31668 31340 31720 31346
rect 31668 31282 31720 31288
rect 31312 30394 31340 31282
rect 31300 30388 31352 30394
rect 31300 30330 31352 30336
rect 31312 29510 31340 30330
rect 31484 30320 31536 30326
rect 31536 30268 31616 30274
rect 31484 30262 31616 30268
rect 31496 30246 31616 30262
rect 31588 30122 31616 30246
rect 31576 30116 31628 30122
rect 31576 30058 31628 30064
rect 31208 29504 31260 29510
rect 31208 29446 31260 29452
rect 31300 29504 31352 29510
rect 31300 29446 31352 29452
rect 31220 29102 31248 29446
rect 31312 29170 31340 29446
rect 31300 29164 31352 29170
rect 31300 29106 31352 29112
rect 31208 29096 31260 29102
rect 31208 29038 31260 29044
rect 30932 28960 30984 28966
rect 30932 28902 30984 28908
rect 30944 28694 30972 28902
rect 31588 28694 31616 30058
rect 31680 30054 31708 31282
rect 31772 30122 31800 31758
rect 32048 31278 32076 32302
rect 32416 31346 32444 33050
rect 32496 32428 32548 32434
rect 32496 32370 32548 32376
rect 32508 31958 32536 32370
rect 32496 31952 32548 31958
rect 32496 31894 32548 31900
rect 32600 31754 32628 34462
rect 32968 34134 32996 37130
rect 33244 35578 33272 37266
rect 34348 36854 34376 37606
rect 34532 37466 34560 37810
rect 34520 37460 34572 37466
rect 34520 37402 34572 37408
rect 34520 37256 34572 37262
rect 34520 37198 34572 37204
rect 34336 36848 34388 36854
rect 34336 36790 34388 36796
rect 34532 35698 34560 37198
rect 34716 37126 34744 39238
rect 34992 38826 35020 39238
rect 35636 39030 35664 40326
rect 35808 39840 35860 39846
rect 35808 39782 35860 39788
rect 35820 39642 35848 39782
rect 35808 39636 35860 39642
rect 35808 39578 35860 39584
rect 35624 39024 35676 39030
rect 35624 38966 35676 38972
rect 34980 38820 35032 38826
rect 34980 38762 35032 38768
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 35912 38350 35940 43046
rect 36268 42696 36320 42702
rect 36268 42638 36320 42644
rect 36280 42226 36308 42638
rect 36452 42628 36504 42634
rect 36452 42570 36504 42576
rect 36464 42362 36492 42570
rect 36452 42356 36504 42362
rect 36452 42298 36504 42304
rect 36268 42220 36320 42226
rect 36268 42162 36320 42168
rect 37096 41676 37148 41682
rect 37096 41618 37148 41624
rect 35992 41132 36044 41138
rect 35992 41074 36044 41080
rect 36004 40050 36032 41074
rect 36084 40928 36136 40934
rect 36084 40870 36136 40876
rect 36268 40928 36320 40934
rect 36268 40870 36320 40876
rect 35992 40044 36044 40050
rect 35992 39986 36044 39992
rect 35440 38344 35492 38350
rect 35440 38286 35492 38292
rect 35900 38344 35952 38350
rect 35900 38286 35952 38292
rect 35348 37800 35400 37806
rect 35348 37742 35400 37748
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34704 37120 34756 37126
rect 34704 37062 34756 37068
rect 34612 36576 34664 36582
rect 34612 36518 34664 36524
rect 34520 35692 34572 35698
rect 34520 35634 34572 35640
rect 33152 35550 33272 35578
rect 33784 35624 33836 35630
rect 33784 35566 33836 35572
rect 32956 34128 33008 34134
rect 32956 34070 33008 34076
rect 33152 33114 33180 35550
rect 33232 35488 33284 35494
rect 33232 35430 33284 35436
rect 33244 35018 33272 35430
rect 33232 35012 33284 35018
rect 33232 34954 33284 34960
rect 33232 34740 33284 34746
rect 33232 34682 33284 34688
rect 33140 33108 33192 33114
rect 33140 33050 33192 33056
rect 33244 32842 33272 34682
rect 33796 34066 33824 35566
rect 34532 34898 34560 35634
rect 34624 35630 34652 36518
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35360 36174 35388 37742
rect 35452 36922 35480 38286
rect 35808 38208 35860 38214
rect 35808 38150 35860 38156
rect 35624 37868 35676 37874
rect 35624 37810 35676 37816
rect 35636 37466 35664 37810
rect 35624 37460 35676 37466
rect 35624 37402 35676 37408
rect 35820 37262 35848 38150
rect 35808 37256 35860 37262
rect 35808 37198 35860 37204
rect 36004 37194 36032 39986
rect 36096 39506 36124 40870
rect 36280 40594 36308 40870
rect 36268 40588 36320 40594
rect 36268 40530 36320 40536
rect 37108 40225 37136 41618
rect 37094 40216 37150 40225
rect 37094 40151 37150 40160
rect 36084 39500 36136 39506
rect 36084 39442 36136 39448
rect 36452 39364 36504 39370
rect 36452 39306 36504 39312
rect 36464 39098 36492 39306
rect 36452 39092 36504 39098
rect 36452 39034 36504 39040
rect 37094 38856 37150 38865
rect 37094 38791 37150 38800
rect 37108 38418 37136 38791
rect 37096 38412 37148 38418
rect 37096 38354 37148 38360
rect 36728 37664 36780 37670
rect 36728 37606 36780 37612
rect 36740 37330 36768 37606
rect 36728 37324 36780 37330
rect 36728 37266 36780 37272
rect 36268 37256 36320 37262
rect 36268 37198 36320 37204
rect 35992 37188 36044 37194
rect 35992 37130 36044 37136
rect 35440 36916 35492 36922
rect 35440 36858 35492 36864
rect 36280 36786 36308 37198
rect 36268 36780 36320 36786
rect 36268 36722 36320 36728
rect 35348 36168 35400 36174
rect 35348 36110 35400 36116
rect 36176 36168 36228 36174
rect 36176 36110 36228 36116
rect 34704 35692 34756 35698
rect 34704 35634 34756 35640
rect 34612 35624 34664 35630
rect 34612 35566 34664 35572
rect 34440 34870 34560 34898
rect 34612 34944 34664 34950
rect 34612 34886 34664 34892
rect 34440 34610 34468 34870
rect 34520 34740 34572 34746
rect 34520 34682 34572 34688
rect 34428 34604 34480 34610
rect 34428 34546 34480 34552
rect 33968 34536 34020 34542
rect 33968 34478 34020 34484
rect 33784 34060 33836 34066
rect 33784 34002 33836 34008
rect 33692 33992 33744 33998
rect 33692 33934 33744 33940
rect 33324 33856 33376 33862
rect 33508 33856 33560 33862
rect 33376 33804 33456 33810
rect 33324 33798 33456 33804
rect 33508 33798 33560 33804
rect 33336 33782 33456 33798
rect 33232 32836 33284 32842
rect 33232 32778 33284 32784
rect 33244 32722 33272 32778
rect 33244 32694 33364 32722
rect 33232 32224 33284 32230
rect 33232 32166 33284 32172
rect 33244 31822 33272 32166
rect 33232 31816 33284 31822
rect 33232 31758 33284 31764
rect 32508 31726 32628 31754
rect 32404 31340 32456 31346
rect 32404 31282 32456 31288
rect 32036 31272 32088 31278
rect 32036 31214 32088 31220
rect 32404 30796 32456 30802
rect 32404 30738 32456 30744
rect 31852 30728 31904 30734
rect 31852 30670 31904 30676
rect 31760 30116 31812 30122
rect 31760 30058 31812 30064
rect 31668 30048 31720 30054
rect 31668 29990 31720 29996
rect 31668 29640 31720 29646
rect 31668 29582 31720 29588
rect 31680 29306 31708 29582
rect 31668 29300 31720 29306
rect 31668 29242 31720 29248
rect 31864 28966 31892 30670
rect 31944 29096 31996 29102
rect 31944 29038 31996 29044
rect 31852 28960 31904 28966
rect 31852 28902 31904 28908
rect 30932 28688 30984 28694
rect 30932 28630 30984 28636
rect 31300 28688 31352 28694
rect 31300 28630 31352 28636
rect 31576 28688 31628 28694
rect 31576 28630 31628 28636
rect 31312 28082 31340 28630
rect 31760 28212 31812 28218
rect 31760 28154 31812 28160
rect 31300 28076 31352 28082
rect 31300 28018 31352 28024
rect 31116 27940 31168 27946
rect 31116 27882 31168 27888
rect 30840 27600 30892 27606
rect 30840 27542 30892 27548
rect 30748 27464 30800 27470
rect 30748 27406 30800 27412
rect 30656 27328 30708 27334
rect 30656 27270 30708 27276
rect 30380 26988 30432 26994
rect 30380 26930 30432 26936
rect 30564 26988 30616 26994
rect 30564 26930 30616 26936
rect 29828 26920 29880 26926
rect 29828 26862 29880 26868
rect 28448 26852 28500 26858
rect 28448 26794 28500 26800
rect 29840 26382 29868 26862
rect 29828 26376 29880 26382
rect 30392 26330 30420 26930
rect 30576 26382 30604 26930
rect 30668 26926 30696 27270
rect 30656 26920 30708 26926
rect 30656 26862 30708 26868
rect 30656 26512 30708 26518
rect 30656 26454 30708 26460
rect 29828 26318 29880 26324
rect 30300 26302 30420 26330
rect 30564 26376 30616 26382
rect 30564 26318 30616 26324
rect 29184 25696 29236 25702
rect 29184 25638 29236 25644
rect 30300 25650 30328 26302
rect 30472 26240 30524 26246
rect 30472 26182 30524 26188
rect 29196 25294 29224 25638
rect 30300 25622 30420 25650
rect 29184 25288 29236 25294
rect 29184 25230 29236 25236
rect 29828 25288 29880 25294
rect 29828 25230 29880 25236
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 28000 23866 28028 24754
rect 29092 24676 29144 24682
rect 29092 24618 29144 24624
rect 28080 24608 28132 24614
rect 28080 24550 28132 24556
rect 28092 24206 28120 24550
rect 28080 24200 28132 24206
rect 28080 24142 28132 24148
rect 28540 24132 28592 24138
rect 28540 24074 28592 24080
rect 28552 23866 28580 24074
rect 27988 23860 28040 23866
rect 27988 23802 28040 23808
rect 28540 23860 28592 23866
rect 28540 23802 28592 23808
rect 27896 23724 27948 23730
rect 27896 23666 27948 23672
rect 27436 23656 27488 23662
rect 27436 23598 27488 23604
rect 27344 23316 27396 23322
rect 27344 23258 27396 23264
rect 27448 23050 27476 23598
rect 27436 23044 27488 23050
rect 27436 22986 27488 22992
rect 26976 22976 27028 22982
rect 26976 22918 27028 22924
rect 26792 22228 26844 22234
rect 26792 22170 26844 22176
rect 26700 22092 26752 22098
rect 26700 22034 26752 22040
rect 26424 21956 26476 21962
rect 26424 21898 26476 21904
rect 26436 21690 26464 21898
rect 26424 21684 26476 21690
rect 26424 21626 26476 21632
rect 26436 21554 26464 21626
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 26424 21548 26476 21554
rect 26424 21490 26476 21496
rect 25056 20466 25084 21490
rect 26516 21344 26568 21350
rect 26516 21286 26568 21292
rect 26528 21146 26556 21286
rect 26516 21140 26568 21146
rect 26516 21082 26568 21088
rect 26712 21010 26740 22034
rect 26804 21486 26832 22170
rect 27804 21888 27856 21894
rect 27804 21830 27856 21836
rect 27816 21554 27844 21830
rect 26976 21548 27028 21554
rect 26976 21490 27028 21496
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 26792 21480 26844 21486
rect 26792 21422 26844 21428
rect 26700 21004 26752 21010
rect 26700 20946 26752 20952
rect 26424 20936 26476 20942
rect 26424 20878 26476 20884
rect 26436 20602 26464 20878
rect 26240 20596 26292 20602
rect 26240 20538 26292 20544
rect 26424 20596 26476 20602
rect 26424 20538 26476 20544
rect 25044 20460 25096 20466
rect 25044 20402 25096 20408
rect 24952 19848 25004 19854
rect 24952 19790 25004 19796
rect 24860 19780 24912 19786
rect 24860 19722 24912 19728
rect 24768 19712 24820 19718
rect 24768 19654 24820 19660
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 24780 19446 24808 19654
rect 24768 19440 24820 19446
rect 24768 19382 24820 19388
rect 24872 18970 24900 19722
rect 25056 19378 25084 20402
rect 26252 20262 26280 20538
rect 26240 20256 26292 20262
rect 26240 20198 26292 20204
rect 26712 19922 26740 20946
rect 26804 20874 26832 21422
rect 26988 21146 27016 21490
rect 26976 21140 27028 21146
rect 26976 21082 27028 21088
rect 26792 20868 26844 20874
rect 26792 20810 26844 20816
rect 26976 20800 27028 20806
rect 26976 20742 27028 20748
rect 27160 20800 27212 20806
rect 27160 20742 27212 20748
rect 26988 20466 27016 20742
rect 27172 20466 27200 20742
rect 27908 20618 27936 23666
rect 28264 23112 28316 23118
rect 28264 23054 28316 23060
rect 28276 22642 28304 23054
rect 28264 22636 28316 22642
rect 28264 22578 28316 22584
rect 28276 22234 28304 22578
rect 28264 22228 28316 22234
rect 28264 22170 28316 22176
rect 27816 20590 27936 20618
rect 26976 20460 27028 20466
rect 26976 20402 27028 20408
rect 27160 20460 27212 20466
rect 27160 20402 27212 20408
rect 26700 19916 26752 19922
rect 26700 19858 26752 19864
rect 26976 19848 27028 19854
rect 26976 19790 27028 19796
rect 26148 19712 26200 19718
rect 26148 19654 26200 19660
rect 26160 19378 26188 19654
rect 26988 19514 27016 19790
rect 26976 19508 27028 19514
rect 26976 19450 27028 19456
rect 27172 19378 27200 20402
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 27632 19514 27660 19790
rect 27816 19718 27844 20590
rect 27896 20460 27948 20466
rect 27896 20402 27948 20408
rect 27804 19712 27856 19718
rect 27804 19654 27856 19660
rect 27620 19508 27672 19514
rect 27620 19450 27672 19456
rect 25044 19372 25096 19378
rect 25044 19314 25096 19320
rect 26148 19372 26200 19378
rect 26148 19314 26200 19320
rect 27160 19372 27212 19378
rect 27160 19314 27212 19320
rect 24860 18964 24912 18970
rect 24860 18906 24912 18912
rect 23296 18624 23348 18630
rect 23296 18566 23348 18572
rect 25056 17746 25084 19314
rect 26608 19168 26660 19174
rect 26608 19110 26660 19116
rect 26620 18766 26648 19110
rect 26608 18760 26660 18766
rect 26608 18702 26660 18708
rect 26792 18760 26844 18766
rect 26792 18702 26844 18708
rect 26804 18630 26832 18702
rect 27172 18630 27200 19314
rect 27252 18828 27304 18834
rect 27252 18770 27304 18776
rect 26424 18624 26476 18630
rect 26424 18566 26476 18572
rect 26792 18624 26844 18630
rect 26792 18566 26844 18572
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 25044 17740 25096 17746
rect 25044 17682 25096 17688
rect 26436 17678 26464 18566
rect 27264 17882 27292 18770
rect 27632 18698 27660 19450
rect 27908 19310 27936 20402
rect 28172 19848 28224 19854
rect 28172 19790 28224 19796
rect 27896 19304 27948 19310
rect 27896 19246 27948 19252
rect 27908 18970 27936 19246
rect 28184 18970 28212 19790
rect 28264 19712 28316 19718
rect 28264 19654 28316 19660
rect 28276 19378 28304 19654
rect 28552 19446 28580 23802
rect 29000 23724 29052 23730
rect 29000 23666 29052 23672
rect 28816 23656 28868 23662
rect 28816 23598 28868 23604
rect 28828 23118 28856 23598
rect 29012 23118 29040 23666
rect 29104 23594 29132 24618
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29748 24206 29776 24550
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 29736 24200 29788 24206
rect 29736 24142 29788 24148
rect 29092 23588 29144 23594
rect 29092 23530 29144 23536
rect 29564 23322 29592 24142
rect 29644 23520 29696 23526
rect 29644 23462 29696 23468
rect 29552 23316 29604 23322
rect 29552 23258 29604 23264
rect 28816 23112 28868 23118
rect 28816 23054 28868 23060
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 28908 23044 28960 23050
rect 28908 22986 28960 22992
rect 28920 22710 28948 22986
rect 28908 22704 28960 22710
rect 28908 22646 28960 22652
rect 29656 22642 29684 23462
rect 29840 23118 29868 25230
rect 30012 24744 30064 24750
rect 30012 24686 30064 24692
rect 30024 24206 30052 24686
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 30012 24200 30064 24206
rect 30012 24142 30064 24148
rect 29932 23730 29960 24142
rect 30024 23730 30052 24142
rect 30104 24132 30156 24138
rect 30104 24074 30156 24080
rect 29920 23724 29972 23730
rect 29920 23666 29972 23672
rect 30012 23724 30064 23730
rect 30012 23666 30064 23672
rect 30116 23594 30144 24074
rect 30196 24064 30248 24070
rect 30196 24006 30248 24012
rect 30392 24018 30420 25622
rect 30484 25158 30512 26182
rect 30668 25906 30696 26454
rect 30656 25900 30708 25906
rect 30656 25842 30708 25848
rect 30472 25152 30524 25158
rect 30472 25094 30524 25100
rect 30484 24614 30512 25094
rect 30472 24608 30524 24614
rect 30472 24550 30524 24556
rect 30760 24206 30788 27406
rect 30852 26994 30880 27542
rect 30840 26988 30892 26994
rect 30840 26930 30892 26936
rect 30932 26920 30984 26926
rect 30932 26862 30984 26868
rect 30944 25838 30972 26862
rect 30932 25832 30984 25838
rect 30932 25774 30984 25780
rect 30748 24200 30800 24206
rect 30748 24142 30800 24148
rect 31024 24132 31076 24138
rect 31024 24074 31076 24080
rect 30748 24064 30800 24070
rect 30208 23730 30236 24006
rect 30392 23990 30512 24018
rect 30748 24006 30800 24012
rect 30196 23724 30248 23730
rect 30196 23666 30248 23672
rect 30104 23588 30156 23594
rect 30104 23530 30156 23536
rect 30116 23254 30144 23530
rect 30104 23248 30156 23254
rect 30104 23190 30156 23196
rect 29828 23112 29880 23118
rect 29828 23054 29880 23060
rect 30104 23112 30156 23118
rect 30104 23054 30156 23060
rect 29736 22976 29788 22982
rect 29736 22918 29788 22924
rect 29748 22642 29776 22918
rect 29644 22636 29696 22642
rect 29644 22578 29696 22584
rect 29736 22636 29788 22642
rect 29736 22578 29788 22584
rect 29828 22568 29880 22574
rect 29828 22510 29880 22516
rect 29552 22500 29604 22506
rect 29552 22442 29604 22448
rect 29092 21344 29144 21350
rect 29092 21286 29144 21292
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 28920 19514 28948 19790
rect 28908 19508 28960 19514
rect 28908 19450 28960 19456
rect 28540 19440 28592 19446
rect 28460 19388 28540 19394
rect 28460 19382 28592 19388
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28460 19366 28580 19382
rect 27896 18964 27948 18970
rect 27896 18906 27948 18912
rect 28172 18964 28224 18970
rect 28172 18906 28224 18912
rect 27620 18692 27672 18698
rect 27620 18634 27672 18640
rect 28460 18290 28488 19366
rect 29104 18698 29132 21286
rect 29564 20398 29592 22442
rect 29840 21146 29868 22510
rect 30116 21554 30144 23054
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 30196 22432 30248 22438
rect 30196 22374 30248 22380
rect 30104 21548 30156 21554
rect 30104 21490 30156 21496
rect 29828 21140 29880 21146
rect 29828 21082 29880 21088
rect 29736 20868 29788 20874
rect 29736 20810 29788 20816
rect 29748 20466 29776 20810
rect 29736 20460 29788 20466
rect 29840 20448 29868 21082
rect 30012 21004 30064 21010
rect 30012 20946 30064 20952
rect 29920 20936 29972 20942
rect 29920 20878 29972 20884
rect 29932 20602 29960 20878
rect 30024 20602 30052 20946
rect 29920 20596 29972 20602
rect 29920 20538 29972 20544
rect 30012 20596 30064 20602
rect 30012 20538 30064 20544
rect 29920 20460 29972 20466
rect 29840 20420 29920 20448
rect 29736 20402 29788 20408
rect 29920 20402 29972 20408
rect 29552 20392 29604 20398
rect 29552 20334 29604 20340
rect 30116 18698 30144 21490
rect 30208 20466 30236 22374
rect 30392 21554 30420 22578
rect 30484 21690 30512 23990
rect 30760 23866 30788 24006
rect 30748 23860 30800 23866
rect 30748 23802 30800 23808
rect 30932 23112 30984 23118
rect 30932 23054 30984 23060
rect 30472 21684 30524 21690
rect 30472 21626 30524 21632
rect 30380 21548 30432 21554
rect 30380 21490 30432 21496
rect 30288 21412 30340 21418
rect 30288 21354 30340 21360
rect 30300 20942 30328 21354
rect 30392 21010 30420 21490
rect 30840 21480 30892 21486
rect 30840 21422 30892 21428
rect 30380 21004 30432 21010
rect 30380 20946 30432 20952
rect 30288 20936 30340 20942
rect 30288 20878 30340 20884
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 30300 20058 30328 20878
rect 30392 20534 30420 20946
rect 30852 20806 30880 21422
rect 30840 20800 30892 20806
rect 30840 20742 30892 20748
rect 30380 20528 30432 20534
rect 30380 20470 30432 20476
rect 30288 20052 30340 20058
rect 30288 19994 30340 20000
rect 30852 19854 30880 20742
rect 30944 20466 30972 23054
rect 31036 22982 31064 24074
rect 31024 22976 31076 22982
rect 31024 22918 31076 22924
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 30944 20058 30972 20402
rect 30932 20052 30984 20058
rect 30932 19994 30984 20000
rect 30840 19848 30892 19854
rect 30840 19790 30892 19796
rect 30852 18766 30880 19790
rect 30840 18760 30892 18766
rect 30840 18702 30892 18708
rect 29092 18692 29144 18698
rect 29092 18634 29144 18640
rect 30104 18692 30156 18698
rect 30104 18634 30156 18640
rect 28540 18624 28592 18630
rect 28540 18566 28592 18572
rect 28552 18290 28580 18566
rect 30116 18426 30144 18634
rect 30104 18420 30156 18426
rect 30104 18362 30156 18368
rect 28448 18284 28500 18290
rect 28448 18226 28500 18232
rect 28540 18284 28592 18290
rect 28540 18226 28592 18232
rect 30852 17882 30880 18702
rect 31128 18222 31156 27882
rect 31392 27396 31444 27402
rect 31392 27338 31444 27344
rect 31404 26586 31432 27338
rect 31392 26580 31444 26586
rect 31392 26522 31444 26528
rect 31772 26466 31800 28154
rect 31680 26438 31800 26466
rect 31680 26382 31708 26438
rect 31668 26376 31720 26382
rect 31668 26318 31720 26324
rect 31484 26240 31536 26246
rect 31484 26182 31536 26188
rect 31496 25838 31524 26182
rect 31484 25832 31536 25838
rect 31484 25774 31536 25780
rect 31772 24818 31800 26438
rect 31852 26036 31904 26042
rect 31852 25978 31904 25984
rect 31864 25906 31892 25978
rect 31852 25900 31904 25906
rect 31852 25842 31904 25848
rect 31760 24812 31812 24818
rect 31760 24754 31812 24760
rect 31772 24274 31800 24754
rect 31760 24268 31812 24274
rect 31760 24210 31812 24216
rect 31208 22976 31260 22982
rect 31208 22918 31260 22924
rect 31220 22642 31248 22918
rect 31208 22636 31260 22642
rect 31208 22578 31260 22584
rect 31484 21548 31536 21554
rect 31484 21490 31536 21496
rect 31208 21412 31260 21418
rect 31208 21354 31260 21360
rect 31220 20942 31248 21354
rect 31392 21344 31444 21350
rect 31392 21286 31444 21292
rect 31404 21010 31432 21286
rect 31496 21010 31524 21490
rect 31956 21146 31984 29038
rect 32036 28620 32088 28626
rect 32036 28562 32088 28568
rect 32048 26790 32076 28562
rect 32036 26784 32088 26790
rect 32036 26726 32088 26732
rect 32048 26382 32076 26726
rect 32128 26444 32180 26450
rect 32128 26386 32180 26392
rect 32036 26376 32088 26382
rect 32036 26318 32088 26324
rect 32140 26042 32168 26386
rect 32128 26036 32180 26042
rect 32128 25978 32180 25984
rect 32220 25832 32272 25838
rect 32220 25774 32272 25780
rect 32232 25498 32260 25774
rect 32220 25492 32272 25498
rect 32220 25434 32272 25440
rect 32036 25288 32088 25294
rect 32036 25230 32088 25236
rect 32048 24954 32076 25230
rect 32036 24948 32088 24954
rect 32036 24890 32088 24896
rect 32312 23792 32364 23798
rect 32312 23734 32364 23740
rect 32128 23044 32180 23050
rect 32128 22986 32180 22992
rect 32140 22778 32168 22986
rect 32128 22772 32180 22778
rect 32128 22714 32180 22720
rect 32128 22024 32180 22030
rect 32128 21966 32180 21972
rect 32220 22024 32272 22030
rect 32220 21966 32272 21972
rect 32140 21690 32168 21966
rect 32128 21684 32180 21690
rect 32128 21626 32180 21632
rect 31944 21140 31996 21146
rect 31944 21082 31996 21088
rect 31392 21004 31444 21010
rect 31392 20946 31444 20952
rect 31484 21004 31536 21010
rect 31484 20946 31536 20952
rect 31208 20936 31260 20942
rect 31208 20878 31260 20884
rect 31852 20800 31904 20806
rect 31852 20742 31904 20748
rect 31668 20528 31720 20534
rect 31668 20470 31720 20476
rect 31680 19854 31708 20470
rect 31760 20324 31812 20330
rect 31760 20266 31812 20272
rect 31668 19848 31720 19854
rect 31668 19790 31720 19796
rect 31772 18834 31800 20266
rect 31760 18828 31812 18834
rect 31760 18770 31812 18776
rect 31864 18766 31892 20742
rect 31852 18760 31904 18766
rect 31852 18702 31904 18708
rect 31300 18624 31352 18630
rect 31300 18566 31352 18572
rect 31576 18624 31628 18630
rect 31576 18566 31628 18572
rect 31312 18290 31340 18566
rect 31588 18290 31616 18566
rect 32232 18426 32260 21966
rect 32324 18698 32352 23734
rect 32312 18692 32364 18698
rect 32312 18634 32364 18640
rect 32220 18420 32272 18426
rect 32220 18362 32272 18368
rect 31300 18284 31352 18290
rect 31300 18226 31352 18232
rect 31576 18284 31628 18290
rect 31576 18226 31628 18232
rect 31116 18216 31168 18222
rect 31116 18158 31168 18164
rect 31208 18080 31260 18086
rect 31208 18022 31260 18028
rect 27252 17876 27304 17882
rect 27252 17818 27304 17824
rect 30840 17876 30892 17882
rect 30840 17818 30892 17824
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 31220 17610 31248 18022
rect 31208 17604 31260 17610
rect 31208 17546 31260 17552
rect 32416 16574 32444 30738
rect 32508 20262 32536 31726
rect 33244 30122 33272 31758
rect 33336 30326 33364 32694
rect 33324 30320 33376 30326
rect 33324 30262 33376 30268
rect 33232 30116 33284 30122
rect 33232 30058 33284 30064
rect 33244 29578 33272 30058
rect 33336 29782 33364 30262
rect 33324 29776 33376 29782
rect 33324 29718 33376 29724
rect 33428 29594 33456 33782
rect 33520 32502 33548 33798
rect 33704 33658 33732 33934
rect 33692 33652 33744 33658
rect 33692 33594 33744 33600
rect 33980 33386 34008 34478
rect 34532 34066 34560 34682
rect 34624 34678 34652 34886
rect 34612 34672 34664 34678
rect 34612 34614 34664 34620
rect 34520 34060 34572 34066
rect 34520 34002 34572 34008
rect 34624 33930 34652 34614
rect 34716 34202 34744 35634
rect 35440 35624 35492 35630
rect 35440 35566 35492 35572
rect 34796 35488 34848 35494
rect 34796 35430 34848 35436
rect 34808 35018 34836 35430
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34796 35012 34848 35018
rect 34796 34954 34848 34960
rect 35452 34610 35480 35566
rect 36188 35086 36216 36110
rect 36360 36100 36412 36106
rect 36360 36042 36412 36048
rect 36372 35834 36400 36042
rect 36360 35828 36412 35834
rect 36360 35770 36412 35776
rect 36544 35692 36596 35698
rect 36544 35634 36596 35640
rect 36556 35290 36584 35634
rect 36544 35284 36596 35290
rect 36544 35226 36596 35232
rect 36360 35148 36412 35154
rect 36360 35090 36412 35096
rect 36176 35080 36228 35086
rect 36176 35022 36228 35028
rect 35808 35012 35860 35018
rect 35808 34954 35860 34960
rect 35440 34604 35492 34610
rect 35440 34546 35492 34552
rect 34796 34400 34848 34406
rect 34796 34342 34848 34348
rect 34704 34196 34756 34202
rect 34704 34138 34756 34144
rect 34612 33924 34664 33930
rect 34612 33866 34664 33872
rect 34808 33522 34836 34342
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 35714 34096 35770 34105
rect 35820 34066 35848 34954
rect 35900 34672 35952 34678
rect 35900 34614 35952 34620
rect 35912 34202 35940 34614
rect 35900 34196 35952 34202
rect 35900 34138 35952 34144
rect 36188 34066 36216 35022
rect 36372 34542 36400 35090
rect 36740 34678 36768 37266
rect 37004 34740 37056 34746
rect 37004 34682 37056 34688
rect 36728 34672 36780 34678
rect 36728 34614 36780 34620
rect 36360 34536 36412 34542
rect 36360 34478 36412 34484
rect 36372 34406 36400 34478
rect 36360 34400 36412 34406
rect 36360 34342 36412 34348
rect 35714 34031 35770 34040
rect 35808 34060 35860 34066
rect 34428 33516 34480 33522
rect 34428 33458 34480 33464
rect 34796 33516 34848 33522
rect 34796 33458 34848 33464
rect 33968 33380 34020 33386
rect 33968 33322 34020 33328
rect 33508 32496 33560 32502
rect 33508 32438 33560 32444
rect 34440 32026 34468 33458
rect 34520 33380 34572 33386
rect 34520 33322 34572 33328
rect 34532 32978 34560 33322
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 34520 32972 34572 32978
rect 34520 32914 34572 32920
rect 35440 32224 35492 32230
rect 35440 32166 35492 32172
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 34428 32020 34480 32026
rect 34428 31962 34480 31968
rect 34060 31272 34112 31278
rect 34060 31214 34112 31220
rect 33784 31136 33836 31142
rect 33784 31078 33836 31084
rect 33692 30048 33744 30054
rect 33692 29990 33744 29996
rect 33232 29572 33284 29578
rect 33232 29514 33284 29520
rect 33336 29566 33456 29594
rect 32864 28416 32916 28422
rect 32864 28358 32916 28364
rect 32772 26784 32824 26790
rect 32772 26726 32824 26732
rect 32680 24064 32732 24070
rect 32680 24006 32732 24012
rect 32692 23526 32720 24006
rect 32680 23520 32732 23526
rect 32680 23462 32732 23468
rect 32692 23118 32720 23462
rect 32680 23112 32732 23118
rect 32680 23054 32732 23060
rect 32588 22636 32640 22642
rect 32588 22578 32640 22584
rect 32600 22234 32628 22578
rect 32588 22228 32640 22234
rect 32588 22170 32640 22176
rect 32588 21480 32640 21486
rect 32588 21422 32640 21428
rect 32600 20942 32628 21422
rect 32588 20936 32640 20942
rect 32588 20878 32640 20884
rect 32496 20256 32548 20262
rect 32496 20198 32548 20204
rect 32692 18290 32720 23054
rect 32784 22642 32812 26726
rect 32876 26382 32904 28358
rect 32956 28076 33008 28082
rect 32956 28018 33008 28024
rect 32968 27606 32996 28018
rect 32956 27600 33008 27606
rect 32956 27542 33008 27548
rect 33336 27418 33364 29566
rect 33416 29504 33468 29510
rect 33416 29446 33468 29452
rect 33428 28558 33456 29446
rect 33704 28626 33732 29990
rect 33796 29714 33824 31078
rect 34072 30258 34100 31214
rect 34440 30326 34468 31962
rect 35348 31952 35400 31958
rect 35348 31894 35400 31900
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34428 30320 34480 30326
rect 34428 30262 34480 30268
rect 34060 30252 34112 30258
rect 34060 30194 34112 30200
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34796 29776 34848 29782
rect 34796 29718 34848 29724
rect 33784 29708 33836 29714
rect 33784 29650 33836 29656
rect 33796 29170 33824 29650
rect 34612 29640 34664 29646
rect 34612 29582 34664 29588
rect 34428 29572 34480 29578
rect 34428 29514 34480 29520
rect 34440 29170 34468 29514
rect 34520 29504 34572 29510
rect 34520 29446 34572 29452
rect 33784 29164 33836 29170
rect 33784 29106 33836 29112
rect 34428 29164 34480 29170
rect 34428 29106 34480 29112
rect 33692 28620 33744 28626
rect 33692 28562 33744 28568
rect 33416 28552 33468 28558
rect 33416 28494 33468 28500
rect 33428 28422 33456 28494
rect 33416 28416 33468 28422
rect 33416 28358 33468 28364
rect 33428 28082 33456 28358
rect 33416 28076 33468 28082
rect 33416 28018 33468 28024
rect 33428 27538 33456 28018
rect 33704 28014 33732 28562
rect 33784 28552 33836 28558
rect 33784 28494 33836 28500
rect 33968 28552 34020 28558
rect 33968 28494 34020 28500
rect 33796 28082 33824 28494
rect 33980 28218 34008 28494
rect 34532 28490 34560 29446
rect 34624 29170 34652 29582
rect 34612 29164 34664 29170
rect 34612 29106 34664 29112
rect 34612 28960 34664 28966
rect 34612 28902 34664 28908
rect 34624 28626 34652 28902
rect 34612 28620 34664 28626
rect 34612 28562 34664 28568
rect 34808 28558 34836 29718
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34796 28552 34848 28558
rect 34796 28494 34848 28500
rect 34520 28484 34572 28490
rect 34520 28426 34572 28432
rect 33968 28212 34020 28218
rect 33968 28154 34020 28160
rect 34532 28082 34560 28426
rect 33784 28076 33836 28082
rect 33784 28018 33836 28024
rect 34520 28076 34572 28082
rect 34520 28018 34572 28024
rect 33692 28008 33744 28014
rect 33692 27950 33744 27956
rect 33508 27940 33560 27946
rect 33508 27882 33560 27888
rect 33416 27532 33468 27538
rect 33416 27474 33468 27480
rect 33520 27470 33548 27882
rect 34060 27872 34112 27878
rect 34060 27814 34112 27820
rect 33508 27464 33560 27470
rect 33336 27390 33456 27418
rect 33508 27406 33560 27412
rect 33324 27328 33376 27334
rect 33324 27270 33376 27276
rect 32956 26580 33008 26586
rect 32956 26522 33008 26528
rect 32864 26376 32916 26382
rect 32864 26318 32916 26324
rect 32876 25294 32904 26318
rect 32864 25288 32916 25294
rect 32864 25230 32916 25236
rect 32968 24818 32996 26522
rect 33336 26450 33364 27270
rect 33324 26444 33376 26450
rect 33324 26386 33376 26392
rect 33048 26376 33100 26382
rect 33048 26318 33100 26324
rect 33060 26042 33088 26318
rect 33232 26308 33284 26314
rect 33232 26250 33284 26256
rect 33244 26042 33272 26250
rect 33048 26036 33100 26042
rect 33048 25978 33100 25984
rect 33232 26036 33284 26042
rect 33232 25978 33284 25984
rect 32956 24812 33008 24818
rect 32956 24754 33008 24760
rect 32968 23798 32996 24754
rect 32956 23792 33008 23798
rect 32956 23734 33008 23740
rect 33060 23610 33088 25978
rect 33428 24410 33456 27390
rect 33508 26784 33560 26790
rect 33508 26726 33560 26732
rect 33520 26382 33548 26726
rect 34072 26382 34100 27814
rect 34808 27402 34836 28494
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34796 27396 34848 27402
rect 34796 27338 34848 27344
rect 34152 26988 34204 26994
rect 34152 26930 34204 26936
rect 34164 26586 34192 26930
rect 34520 26784 34572 26790
rect 34520 26726 34572 26732
rect 34152 26580 34204 26586
rect 34152 26522 34204 26528
rect 34532 26450 34560 26726
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 35360 26625 35388 31894
rect 35452 31414 35480 32166
rect 35440 31408 35492 31414
rect 35440 31350 35492 31356
rect 35440 30048 35492 30054
rect 35440 29990 35492 29996
rect 35452 29714 35480 29990
rect 35440 29708 35492 29714
rect 35440 29650 35492 29656
rect 35624 29164 35676 29170
rect 35624 29106 35676 29112
rect 35636 27826 35664 29106
rect 35728 28014 35756 34031
rect 35808 34002 35860 34008
rect 36176 34060 36228 34066
rect 36176 34002 36228 34008
rect 35820 32978 35848 34002
rect 36188 32978 36216 34002
rect 37016 33930 37044 34682
rect 36268 33924 36320 33930
rect 36268 33866 36320 33872
rect 37004 33924 37056 33930
rect 37004 33866 37056 33872
rect 36280 33590 36308 33866
rect 36268 33584 36320 33590
rect 36268 33526 36320 33532
rect 35808 32972 35860 32978
rect 35808 32914 35860 32920
rect 36176 32972 36228 32978
rect 36176 32914 36228 32920
rect 35820 32502 35848 32914
rect 35808 32496 35860 32502
rect 35808 32438 35860 32444
rect 36280 32434 36308 33526
rect 36452 33312 36504 33318
rect 36452 33254 36504 33260
rect 36464 32910 36492 33254
rect 36452 32904 36504 32910
rect 36452 32846 36504 32852
rect 36268 32428 36320 32434
rect 36268 32370 36320 32376
rect 37200 31754 37228 47398
rect 37384 46034 37412 49200
rect 37740 47048 37792 47054
rect 37740 46990 37792 46996
rect 37372 46028 37424 46034
rect 37372 45970 37424 45976
rect 37372 45892 37424 45898
rect 37372 45834 37424 45840
rect 37384 45558 37412 45834
rect 37372 45552 37424 45558
rect 37372 45494 37424 45500
rect 37280 45484 37332 45490
rect 37280 45426 37332 45432
rect 37292 37874 37320 45426
rect 37372 45076 37424 45082
rect 37372 45018 37424 45024
rect 37384 44402 37412 45018
rect 37752 45014 37780 46990
rect 38016 46572 38068 46578
rect 38016 46514 38068 46520
rect 38028 45830 38056 46514
rect 38016 45824 38068 45830
rect 38016 45766 38068 45772
rect 37924 45280 37976 45286
rect 37924 45222 37976 45228
rect 37740 45008 37792 45014
rect 37740 44950 37792 44956
rect 37936 44946 37964 45222
rect 37924 44940 37976 44946
rect 37924 44882 37976 44888
rect 37372 44396 37424 44402
rect 37372 44338 37424 44344
rect 37372 44260 37424 44266
rect 37372 44202 37424 44208
rect 37384 42226 37412 44202
rect 37464 43716 37516 43722
rect 37464 43658 37516 43664
rect 37476 43450 37504 43658
rect 37464 43444 37516 43450
rect 37464 43386 37516 43392
rect 37832 43308 37884 43314
rect 37832 43250 37884 43256
rect 37844 42906 37872 43250
rect 37832 42900 37884 42906
rect 37832 42842 37884 42848
rect 37372 42220 37424 42226
rect 37372 42162 37424 42168
rect 37384 40610 37412 42162
rect 37464 41540 37516 41546
rect 37464 41482 37516 41488
rect 37476 41274 37504 41482
rect 37464 41268 37516 41274
rect 37464 41210 37516 41216
rect 37384 40582 37504 40610
rect 37372 40452 37424 40458
rect 37372 40394 37424 40400
rect 37384 40050 37412 40394
rect 37372 40044 37424 40050
rect 37372 39986 37424 39992
rect 37476 38962 37504 40582
rect 37464 38956 37516 38962
rect 37464 38898 37516 38904
rect 37464 38276 37516 38282
rect 37464 38218 37516 38224
rect 37476 38010 37504 38218
rect 37464 38004 37516 38010
rect 37464 37946 37516 37952
rect 37280 37868 37332 37874
rect 37280 37810 37332 37816
rect 37464 37188 37516 37194
rect 37464 37130 37516 37136
rect 37476 36922 37504 37130
rect 37464 36916 37516 36922
rect 37464 36858 37516 36864
rect 37372 36780 37424 36786
rect 37372 36722 37424 36728
rect 37384 36378 37412 36722
rect 37372 36372 37424 36378
rect 37372 36314 37424 36320
rect 37464 36032 37516 36038
rect 37464 35974 37516 35980
rect 37476 35086 37504 35974
rect 37464 35080 37516 35086
rect 37464 35022 37516 35028
rect 37476 33998 37504 35022
rect 37556 34944 37608 34950
rect 37556 34886 37608 34892
rect 37568 34610 37596 34886
rect 37556 34604 37608 34610
rect 37556 34546 37608 34552
rect 37740 34196 37792 34202
rect 37740 34138 37792 34144
rect 37464 33992 37516 33998
rect 37464 33934 37516 33940
rect 37280 33516 37332 33522
rect 37280 33458 37332 33464
rect 37292 32570 37320 33458
rect 37476 33318 37504 33934
rect 37556 33856 37608 33862
rect 37556 33798 37608 33804
rect 37568 33522 37596 33798
rect 37752 33522 37780 34138
rect 37556 33516 37608 33522
rect 37556 33458 37608 33464
rect 37740 33516 37792 33522
rect 37740 33458 37792 33464
rect 37464 33312 37516 33318
rect 37464 33254 37516 33260
rect 37568 33114 37596 33458
rect 37556 33108 37608 33114
rect 37556 33050 37608 33056
rect 37280 32564 37332 32570
rect 37280 32506 37332 32512
rect 37752 32434 37780 33458
rect 37740 32428 37792 32434
rect 37740 32370 37792 32376
rect 37464 31884 37516 31890
rect 37464 31826 37516 31832
rect 37108 31726 37228 31754
rect 36268 30048 36320 30054
rect 36268 29990 36320 29996
rect 36280 29714 36308 29990
rect 36268 29708 36320 29714
rect 36268 29650 36320 29656
rect 35806 29336 35862 29345
rect 35806 29271 35862 29280
rect 35820 29238 35848 29271
rect 35808 29232 35860 29238
rect 35808 29174 35860 29180
rect 35808 28960 35860 28966
rect 35808 28902 35860 28908
rect 36728 28960 36780 28966
rect 36728 28902 36780 28908
rect 35820 28626 35848 28902
rect 35808 28620 35860 28626
rect 35808 28562 35860 28568
rect 36084 28416 36136 28422
rect 36084 28358 36136 28364
rect 35716 28008 35768 28014
rect 35716 27950 35768 27956
rect 35636 27798 35756 27826
rect 35728 27062 35756 27798
rect 35716 27056 35768 27062
rect 35716 26998 35768 27004
rect 35624 26784 35676 26790
rect 35624 26726 35676 26732
rect 35346 26616 35402 26625
rect 35346 26551 35402 26560
rect 34520 26444 34572 26450
rect 34520 26386 34572 26392
rect 34704 26444 34756 26450
rect 34704 26386 34756 26392
rect 35348 26444 35400 26450
rect 35348 26386 35400 26392
rect 33508 26376 33560 26382
rect 33508 26318 33560 26324
rect 34060 26376 34112 26382
rect 34060 26318 34112 26324
rect 33784 25900 33836 25906
rect 33784 25842 33836 25848
rect 33600 24676 33652 24682
rect 33600 24618 33652 24624
rect 33140 24404 33192 24410
rect 33140 24346 33192 24352
rect 33416 24404 33468 24410
rect 33416 24346 33468 24352
rect 32876 23594 33088 23610
rect 32864 23588 33088 23594
rect 32916 23582 33088 23588
rect 32864 23530 32916 23536
rect 32876 22710 32904 23530
rect 32864 22704 32916 22710
rect 32864 22646 32916 22652
rect 32772 22636 32824 22642
rect 32772 22578 32824 22584
rect 33048 21548 33100 21554
rect 33048 21490 33100 21496
rect 32772 21412 32824 21418
rect 32772 21354 32824 21360
rect 32784 20942 32812 21354
rect 32772 20936 32824 20942
rect 32772 20878 32824 20884
rect 33060 20874 33088 21490
rect 33152 21350 33180 24346
rect 33428 24206 33456 24346
rect 33612 24206 33640 24618
rect 33692 24608 33744 24614
rect 33692 24550 33744 24556
rect 33704 24274 33732 24550
rect 33796 24274 33824 25842
rect 33968 24744 34020 24750
rect 33968 24686 34020 24692
rect 33692 24268 33744 24274
rect 33692 24210 33744 24216
rect 33784 24268 33836 24274
rect 33784 24210 33836 24216
rect 33416 24200 33468 24206
rect 33416 24142 33468 24148
rect 33600 24200 33652 24206
rect 33600 24142 33652 24148
rect 33600 23724 33652 23730
rect 33600 23666 33652 23672
rect 33612 23118 33640 23666
rect 33796 23254 33824 24210
rect 33980 23662 34008 24686
rect 34072 23730 34100 26318
rect 34520 26240 34572 26246
rect 34520 26182 34572 26188
rect 34532 25906 34560 26182
rect 34520 25900 34572 25906
rect 34520 25842 34572 25848
rect 34532 25430 34560 25842
rect 34716 25702 34744 26386
rect 34980 26376 35032 26382
rect 34980 26318 35032 26324
rect 34992 26042 35020 26318
rect 34980 26036 35032 26042
rect 34980 25978 35032 25984
rect 35360 25906 35388 26386
rect 34796 25900 34848 25906
rect 34796 25842 34848 25848
rect 34980 25900 35032 25906
rect 35348 25900 35400 25906
rect 35032 25860 35348 25888
rect 34980 25842 35032 25848
rect 35348 25842 35400 25848
rect 34704 25696 34756 25702
rect 34704 25638 34756 25644
rect 34520 25424 34572 25430
rect 34520 25366 34572 25372
rect 34152 24812 34204 24818
rect 34152 24754 34204 24760
rect 34164 24614 34192 24754
rect 34520 24744 34572 24750
rect 34520 24686 34572 24692
rect 34152 24608 34204 24614
rect 34152 24550 34204 24556
rect 34532 23866 34560 24686
rect 34716 24614 34744 25638
rect 34808 25362 34836 25842
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34796 25356 34848 25362
rect 34796 25298 34848 25304
rect 34888 25288 34940 25294
rect 34888 25230 34940 25236
rect 35348 25288 35400 25294
rect 35348 25230 35400 25236
rect 34796 25152 34848 25158
rect 34796 25094 34848 25100
rect 34704 24608 34756 24614
rect 34704 24550 34756 24556
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 34060 23724 34112 23730
rect 34060 23666 34112 23672
rect 33968 23656 34020 23662
rect 33968 23598 34020 23604
rect 33784 23248 33836 23254
rect 33704 23196 33784 23202
rect 33704 23190 33836 23196
rect 33704 23174 33824 23190
rect 33600 23112 33652 23118
rect 33600 23054 33652 23060
rect 33612 22778 33640 23054
rect 33600 22772 33652 22778
rect 33600 22714 33652 22720
rect 33704 22030 33732 23174
rect 33980 22094 34008 23598
rect 34244 22568 34296 22574
rect 34244 22510 34296 22516
rect 34520 22568 34572 22574
rect 34520 22510 34572 22516
rect 34256 22234 34284 22510
rect 34244 22228 34296 22234
rect 34244 22170 34296 22176
rect 33796 22066 34008 22094
rect 34428 22092 34480 22098
rect 33692 22024 33744 22030
rect 33692 21966 33744 21972
rect 33796 21672 33824 22066
rect 34428 22034 34480 22040
rect 33704 21644 33824 21672
rect 33324 21548 33376 21554
rect 33324 21490 33376 21496
rect 33140 21344 33192 21350
rect 33140 21286 33192 21292
rect 33048 20868 33100 20874
rect 33048 20810 33100 20816
rect 33060 20602 33088 20810
rect 33048 20596 33100 20602
rect 33048 20538 33100 20544
rect 33140 20528 33192 20534
rect 33140 20470 33192 20476
rect 33152 20398 33180 20470
rect 33140 20392 33192 20398
rect 33140 20334 33192 20340
rect 33152 19378 33180 20334
rect 33336 20058 33364 21490
rect 33704 20806 33732 21644
rect 34440 21554 34468 22034
rect 34532 21690 34560 22510
rect 34612 22500 34664 22506
rect 34612 22442 34664 22448
rect 34520 21684 34572 21690
rect 34520 21626 34572 21632
rect 34428 21548 34480 21554
rect 34428 21490 34480 21496
rect 34440 21010 34468 21490
rect 34532 21010 34560 21626
rect 34428 21004 34480 21010
rect 34428 20946 34480 20952
rect 34520 21004 34572 21010
rect 34520 20946 34572 20952
rect 34624 20942 34652 22442
rect 34808 22030 34836 25094
rect 34900 24954 34928 25230
rect 34888 24948 34940 24954
rect 34888 24890 34940 24896
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 35360 24410 35388 25230
rect 35636 24410 35664 26726
rect 35348 24404 35400 24410
rect 35348 24346 35400 24352
rect 35624 24404 35676 24410
rect 35624 24346 35676 24352
rect 35440 24200 35492 24206
rect 35440 24142 35492 24148
rect 35348 23724 35400 23730
rect 35348 23666 35400 23672
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 34808 21554 34836 21966
rect 35360 21570 35388 23666
rect 35452 23118 35480 24142
rect 35532 24064 35584 24070
rect 35532 24006 35584 24012
rect 35544 23798 35572 24006
rect 35636 23866 35664 24346
rect 35624 23860 35676 23866
rect 35624 23802 35676 23808
rect 35532 23792 35584 23798
rect 35532 23734 35584 23740
rect 35440 23112 35492 23118
rect 35440 23054 35492 23060
rect 35532 22976 35584 22982
rect 35532 22918 35584 22924
rect 35544 22098 35572 22918
rect 35624 22432 35676 22438
rect 35624 22374 35676 22380
rect 35532 22092 35584 22098
rect 35532 22034 35584 22040
rect 35176 21554 35388 21570
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 35164 21548 35388 21554
rect 35216 21542 35388 21548
rect 35164 21490 35216 21496
rect 33784 20936 33836 20942
rect 33784 20878 33836 20884
rect 34060 20936 34112 20942
rect 34060 20878 34112 20884
rect 34612 20936 34664 20942
rect 34612 20878 34664 20884
rect 33692 20800 33744 20806
rect 33692 20742 33744 20748
rect 33704 20602 33732 20742
rect 33692 20596 33744 20602
rect 33692 20538 33744 20544
rect 33704 20330 33732 20538
rect 33692 20324 33744 20330
rect 33692 20266 33744 20272
rect 33324 20052 33376 20058
rect 33324 19994 33376 20000
rect 33704 19854 33732 20266
rect 33692 19848 33744 19854
rect 33692 19790 33744 19796
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 33152 18834 33180 19314
rect 33796 19310 33824 20878
rect 34072 20602 34100 20878
rect 34060 20596 34112 20602
rect 34060 20538 34112 20544
rect 34336 20460 34388 20466
rect 34336 20402 34388 20408
rect 34244 19372 34296 19378
rect 34244 19314 34296 19320
rect 33784 19304 33836 19310
rect 33784 19246 33836 19252
rect 33140 18828 33192 18834
rect 33140 18770 33192 18776
rect 33796 18766 33824 19246
rect 33784 18760 33836 18766
rect 33784 18702 33836 18708
rect 32956 18624 33008 18630
rect 32956 18566 33008 18572
rect 32680 18284 32732 18290
rect 32680 18226 32732 18232
rect 32692 17746 32720 18226
rect 32772 18216 32824 18222
rect 32772 18158 32824 18164
rect 32784 17746 32812 18158
rect 32968 17882 32996 18566
rect 34256 18426 34284 19314
rect 34348 19310 34376 20402
rect 34624 20330 34652 20878
rect 34808 20874 34836 21490
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34796 20868 34848 20874
rect 34796 20810 34848 20816
rect 35348 20800 35400 20806
rect 35348 20742 35400 20748
rect 34612 20324 34664 20330
rect 34612 20266 34664 20272
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34336 19304 34388 19310
rect 34336 19246 34388 19252
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 35360 18834 35388 20742
rect 35544 20466 35572 22034
rect 35636 21554 35664 22374
rect 35624 21548 35676 21554
rect 35624 21490 35676 21496
rect 35532 20460 35584 20466
rect 35532 20402 35584 20408
rect 35348 18828 35400 18834
rect 35348 18770 35400 18776
rect 34704 18624 34756 18630
rect 34704 18566 34756 18572
rect 33140 18420 33192 18426
rect 33140 18362 33192 18368
rect 34244 18420 34296 18426
rect 34244 18362 34296 18368
rect 32956 17876 33008 17882
rect 32956 17818 33008 17824
rect 32680 17740 32732 17746
rect 32680 17682 32732 17688
rect 32772 17740 32824 17746
rect 32772 17682 32824 17688
rect 33152 17678 33180 18362
rect 33232 18284 33284 18290
rect 33232 18226 33284 18232
rect 33244 17814 33272 18226
rect 33232 17808 33284 17814
rect 33232 17750 33284 17756
rect 34716 17678 34744 18566
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 33140 17672 33192 17678
rect 33140 17614 33192 17620
rect 34704 17672 34756 17678
rect 34704 17614 34756 17620
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 32416 16546 32628 16574
rect 24400 4616 24452 4622
rect 24400 4558 24452 4564
rect 23664 4208 23716 4214
rect 23664 4150 23716 4156
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 22204 2854 22232 4082
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 23572 4072 23624 4078
rect 23572 4014 23624 4020
rect 22572 3670 22600 4014
rect 23018 3768 23074 3777
rect 23018 3703 23074 3712
rect 22560 3664 22612 3670
rect 22560 3606 22612 3612
rect 23032 3534 23060 3703
rect 23584 3670 23612 4014
rect 23572 3664 23624 3670
rect 23572 3606 23624 3612
rect 23676 3534 23704 4150
rect 23848 4072 23900 4078
rect 23848 4014 23900 4020
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23664 3528 23716 3534
rect 23664 3470 23716 3476
rect 22192 2848 22244 2854
rect 22192 2790 22244 2796
rect 21732 2644 21784 2650
rect 21732 2586 21784 2592
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 21284 800 21312 2382
rect 22572 800 22600 3470
rect 23860 800 23888 4014
rect 24412 3602 24440 4558
rect 32220 4140 32272 4146
rect 32220 4082 32272 4088
rect 24584 3936 24636 3942
rect 24584 3878 24636 3884
rect 24596 3602 24624 3878
rect 32232 3602 32260 4082
rect 32496 4072 32548 4078
rect 32496 4014 32548 4020
rect 32508 3738 32536 4014
rect 32496 3732 32548 3738
rect 32496 3674 32548 3680
rect 24400 3596 24452 3602
rect 24400 3538 24452 3544
rect 24584 3596 24636 3602
rect 24584 3538 24636 3544
rect 32220 3596 32272 3602
rect 32220 3538 32272 3544
rect 32600 3534 32628 16546
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 35728 6914 35756 26998
rect 36096 26450 36124 28358
rect 36740 28082 36768 28902
rect 37108 28626 37136 31726
rect 37476 31482 37504 31826
rect 37464 31476 37516 31482
rect 37464 31418 37516 31424
rect 37556 31340 37608 31346
rect 37556 31282 37608 31288
rect 37568 31142 37596 31282
rect 37752 31210 37780 32370
rect 37740 31204 37792 31210
rect 37740 31146 37792 31152
rect 37556 31136 37608 31142
rect 37556 31078 37608 31084
rect 37188 30796 37240 30802
rect 37188 30738 37240 30744
rect 37280 30796 37332 30802
rect 37280 30738 37332 30744
rect 37200 30705 37228 30738
rect 37186 30696 37242 30705
rect 37186 30631 37242 30640
rect 37292 30258 37320 30738
rect 37280 30252 37332 30258
rect 37280 30194 37332 30200
rect 37464 30252 37516 30258
rect 37464 30194 37516 30200
rect 37292 29170 37320 30194
rect 37372 29572 37424 29578
rect 37372 29514 37424 29520
rect 37384 29306 37412 29514
rect 37372 29300 37424 29306
rect 37372 29242 37424 29248
rect 37476 29186 37504 30194
rect 37280 29164 37332 29170
rect 37280 29106 37332 29112
rect 37384 29158 37504 29186
rect 37096 28620 37148 28626
rect 37096 28562 37148 28568
rect 36728 28076 36780 28082
rect 36728 28018 36780 28024
rect 37186 27976 37242 27985
rect 37186 27911 37242 27920
rect 37200 27538 37228 27911
rect 37188 27532 37240 27538
rect 37188 27474 37240 27480
rect 36176 27056 36228 27062
rect 36176 26998 36228 27004
rect 36084 26444 36136 26450
rect 36084 26386 36136 26392
rect 35900 24812 35952 24818
rect 35900 24754 35952 24760
rect 35912 24206 35940 24754
rect 36096 24750 36124 26386
rect 36188 26382 36216 26998
rect 37384 26994 37412 29158
rect 37568 29050 37596 31078
rect 37476 29022 37596 29050
rect 37372 26988 37424 26994
rect 37372 26930 37424 26936
rect 37384 26382 37412 26930
rect 37476 26926 37504 29022
rect 37556 28076 37608 28082
rect 37556 28018 37608 28024
rect 37568 27334 37596 28018
rect 37556 27328 37608 27334
rect 37556 27270 37608 27276
rect 37464 26920 37516 26926
rect 37464 26862 37516 26868
rect 36176 26376 36228 26382
rect 36176 26318 36228 26324
rect 37372 26376 37424 26382
rect 37372 26318 37424 26324
rect 37464 26308 37516 26314
rect 37464 26250 37516 26256
rect 37186 25936 37242 25945
rect 37186 25871 37242 25880
rect 36544 25696 36596 25702
rect 36544 25638 36596 25644
rect 36084 24744 36136 24750
rect 36084 24686 36136 24692
rect 36096 24274 36124 24686
rect 36556 24274 36584 25638
rect 37200 25362 37228 25871
rect 37188 25356 37240 25362
rect 37188 25298 37240 25304
rect 36084 24268 36136 24274
rect 36084 24210 36136 24216
rect 36544 24268 36596 24274
rect 36544 24210 36596 24216
rect 35900 24200 35952 24206
rect 35900 24142 35952 24148
rect 35912 23866 35940 24142
rect 37476 24138 37504 26250
rect 37464 24132 37516 24138
rect 37464 24074 37516 24080
rect 37186 23896 37242 23905
rect 35900 23860 35952 23866
rect 37186 23831 37242 23840
rect 35900 23802 35952 23808
rect 37200 23186 37228 23831
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 37188 23180 37240 23186
rect 37188 23122 37240 23128
rect 36268 22636 36320 22642
rect 36268 22578 36320 22584
rect 36280 22030 36308 22578
rect 37188 22092 37240 22098
rect 37188 22034 37240 22040
rect 36268 22024 36320 22030
rect 36268 21966 36320 21972
rect 36280 21690 36308 21966
rect 37200 21865 37228 22034
rect 37186 21856 37242 21865
rect 37186 21791 37242 21800
rect 36268 21684 36320 21690
rect 36268 21626 36320 21632
rect 36268 20936 36320 20942
rect 36268 20878 36320 20884
rect 36280 20466 36308 20878
rect 37186 20496 37242 20505
rect 36268 20460 36320 20466
rect 37186 20431 37242 20440
rect 36268 20402 36320 20408
rect 37200 19922 37228 20431
rect 37188 19916 37240 19922
rect 37188 19858 37240 19864
rect 36268 18760 36320 18766
rect 36268 18702 36320 18708
rect 36280 18290 36308 18702
rect 36452 18692 36504 18698
rect 36452 18634 36504 18640
rect 36464 18426 36492 18634
rect 36452 18420 36504 18426
rect 36452 18362 36504 18368
rect 36268 18284 36320 18290
rect 36268 18226 36320 18232
rect 36084 18080 36136 18086
rect 36084 18022 36136 18028
rect 36096 17746 36124 18022
rect 36084 17740 36136 17746
rect 36084 17682 36136 17688
rect 36452 17604 36504 17610
rect 36452 17546 36504 17552
rect 36464 17338 36492 17546
rect 36452 17332 36504 17338
rect 36452 17274 36504 17280
rect 36268 16992 36320 16998
rect 36268 16934 36320 16940
rect 36280 16658 36308 16934
rect 36268 16652 36320 16658
rect 36268 16594 36320 16600
rect 36452 16516 36504 16522
rect 36452 16458 36504 16464
rect 36464 16250 36492 16458
rect 36452 16244 36504 16250
rect 36452 16186 36504 16192
rect 36268 15904 36320 15910
rect 36268 15846 36320 15852
rect 36280 15570 36308 15846
rect 36268 15564 36320 15570
rect 36268 15506 36320 15512
rect 36452 15428 36504 15434
rect 36452 15370 36504 15376
rect 36464 15162 36492 15370
rect 36452 15156 36504 15162
rect 36452 15098 36504 15104
rect 36360 15020 36412 15026
rect 36360 14962 36412 14968
rect 36268 10056 36320 10062
rect 36268 9998 36320 10004
rect 36280 9586 36308 9998
rect 36268 9580 36320 9586
rect 36268 9522 36320 9528
rect 35636 6886 35756 6914
rect 36372 6914 36400 14962
rect 37186 11656 37242 11665
rect 37186 11591 37242 11600
rect 37200 11218 37228 11591
rect 37188 11212 37240 11218
rect 37188 11154 37240 11160
rect 36452 10464 36504 10470
rect 36452 10406 36504 10412
rect 36464 10130 36492 10406
rect 36452 10124 36504 10130
rect 36452 10066 36504 10072
rect 37186 9616 37242 9625
rect 37186 9551 37242 9560
rect 37200 9042 37228 9551
rect 37188 9036 37240 9042
rect 37188 8978 37240 8984
rect 37186 7576 37242 7585
rect 37186 7511 37242 7520
rect 36372 6886 36492 6914
rect 35348 6248 35400 6254
rect 35348 6190 35400 6196
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 33416 5704 33468 5710
rect 33416 5646 33468 5652
rect 34520 5704 34572 5710
rect 34520 5646 34572 5652
rect 33428 5234 33456 5646
rect 32680 5228 32732 5234
rect 32680 5170 32732 5176
rect 33416 5228 33468 5234
rect 33416 5170 33468 5176
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 32588 3528 32640 3534
rect 32588 3470 32640 3476
rect 24136 3398 24164 3470
rect 27804 3460 27856 3466
rect 27804 3402 27856 3408
rect 24032 3392 24084 3398
rect 24032 3334 24084 3340
rect 24124 3392 24176 3398
rect 24124 3334 24176 3340
rect 24044 3126 24072 3334
rect 24032 3120 24084 3126
rect 24032 3062 24084 3068
rect 27816 3058 27844 3402
rect 27988 3392 28040 3398
rect 27988 3334 28040 3340
rect 28000 3126 28028 3334
rect 27988 3120 28040 3126
rect 27988 3062 28040 3068
rect 27804 3052 27856 3058
rect 27804 2994 27856 3000
rect 24492 2984 24544 2990
rect 24492 2926 24544 2932
rect 28356 2984 28408 2990
rect 28356 2926 28408 2932
rect 24504 800 24532 2926
rect 28368 800 28396 2926
rect 32600 2922 32628 3470
rect 32588 2916 32640 2922
rect 32588 2858 32640 2864
rect 32692 2854 32720 5170
rect 33968 5092 34020 5098
rect 33968 5034 34020 5040
rect 33980 4690 34008 5034
rect 34532 4690 34560 5646
rect 35254 5536 35310 5545
rect 35254 5471 35310 5480
rect 35268 5302 35296 5471
rect 35256 5296 35308 5302
rect 35256 5238 35308 5244
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34612 4752 34664 4758
rect 34612 4694 34664 4700
rect 33968 4684 34020 4690
rect 33968 4626 34020 4632
rect 34520 4684 34572 4690
rect 34520 4626 34572 4632
rect 34624 4185 34652 4694
rect 34610 4176 34666 4185
rect 34610 4111 34666 4120
rect 34152 4072 34204 4078
rect 34980 4072 35032 4078
rect 34152 4014 34204 4020
rect 34808 4020 34980 4026
rect 34808 4014 35032 4020
rect 34164 3738 34192 4014
rect 34808 3998 35020 4014
rect 34808 3738 34836 3998
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 34152 3732 34204 3738
rect 34152 3674 34204 3680
rect 34796 3732 34848 3738
rect 34796 3674 34848 3680
rect 33232 3528 33284 3534
rect 33232 3470 33284 3476
rect 33244 3058 33272 3470
rect 33416 3392 33468 3398
rect 33416 3334 33468 3340
rect 33428 3126 33456 3334
rect 35360 3194 35388 6190
rect 35532 5568 35584 5574
rect 35532 5510 35584 5516
rect 35544 4690 35572 5510
rect 35532 4684 35584 4690
rect 35532 4626 35584 4632
rect 35440 4072 35492 4078
rect 35440 4014 35492 4020
rect 35348 3188 35400 3194
rect 35348 3130 35400 3136
rect 33416 3120 33468 3126
rect 33416 3062 33468 3068
rect 33232 3052 33284 3058
rect 33232 2994 33284 3000
rect 32680 2848 32732 2854
rect 32680 2790 32732 2796
rect 33692 2848 33744 2854
rect 35348 2848 35400 2854
rect 33692 2790 33744 2796
rect 35346 2816 35348 2825
rect 35400 2816 35402 2825
rect 33704 2514 33732 2790
rect 34934 2748 35242 2768
rect 35346 2751 35402 2760
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 33692 2508 33744 2514
rect 33692 2450 33744 2456
rect 35452 800 35480 4014
rect 35636 3534 35664 6886
rect 36464 5710 36492 6886
rect 37200 6866 37228 7511
rect 37188 6860 37240 6866
rect 37188 6802 37240 6808
rect 36544 6248 36596 6254
rect 36544 6190 36596 6196
rect 37186 6216 37242 6225
rect 36452 5704 36504 5710
rect 36452 5646 36504 5652
rect 36556 5370 36584 6190
rect 37186 6151 37242 6160
rect 37200 5778 37228 6151
rect 37188 5772 37240 5778
rect 37188 5714 37240 5720
rect 36544 5364 36596 5370
rect 36544 5306 36596 5312
rect 36084 4684 36136 4690
rect 36084 4626 36136 4632
rect 35624 3528 35676 3534
rect 35624 3470 35676 3476
rect 35808 3460 35860 3466
rect 35808 3402 35860 3408
rect 35716 3392 35768 3398
rect 35716 3334 35768 3340
rect 35532 2984 35584 2990
rect 35532 2926 35584 2932
rect 35544 1465 35572 2926
rect 35728 2378 35756 3334
rect 35716 2372 35768 2378
rect 35716 2314 35768 2320
rect 35530 1456 35586 1465
rect 35530 1391 35586 1400
rect -10 0 102 800
rect 634 0 746 800
rect 1278 0 1390 800
rect 1922 0 2034 800
rect 3210 0 3322 800
rect 3854 0 3966 800
rect 4498 0 4610 800
rect 5142 0 5254 800
rect 6430 0 6542 800
rect 7074 0 7186 800
rect 7718 0 7830 800
rect 9006 0 9118 800
rect 9650 0 9762 800
rect 10294 0 10406 800
rect 10938 0 11050 800
rect 12226 0 12338 800
rect 12870 0 12982 800
rect 13514 0 13626 800
rect 14802 0 14914 800
rect 15446 0 15558 800
rect 16090 0 16202 800
rect 16734 0 16846 800
rect 18022 0 18134 800
rect 18666 0 18778 800
rect 19310 0 19422 800
rect 20598 0 20710 800
rect 21242 0 21354 800
rect 21886 0 21998 800
rect 22530 0 22642 800
rect 23818 0 23930 800
rect 24462 0 24574 800
rect 25106 0 25218 800
rect 26394 0 26506 800
rect 27038 0 27150 800
rect 27682 0 27794 800
rect 28326 0 28438 800
rect 29614 0 29726 800
rect 30258 0 30370 800
rect 30902 0 31014 800
rect 32190 0 32302 800
rect 32834 0 32946 800
rect 33478 0 33590 800
rect 34122 0 34234 800
rect 35410 0 35522 800
rect 35820 785 35848 3402
rect 35992 2848 36044 2854
rect 35992 2790 36044 2796
rect 36004 2514 36032 2790
rect 35992 2508 36044 2514
rect 35992 2450 36044 2456
rect 36096 800 36124 4626
rect 37292 4146 37320 23666
rect 37464 21956 37516 21962
rect 37464 21898 37516 21904
rect 37476 21690 37504 21898
rect 37464 21684 37516 21690
rect 37464 21626 37516 21632
rect 37464 18284 37516 18290
rect 37464 18226 37516 18232
rect 37476 17202 37504 18226
rect 37464 17196 37516 17202
rect 37464 17138 37516 17144
rect 37464 16108 37516 16114
rect 37464 16050 37516 16056
rect 37372 11756 37424 11762
rect 37372 11698 37424 11704
rect 37384 6914 37412 11698
rect 37476 9586 37504 16050
rect 37568 10674 37596 27270
rect 37844 27146 37872 42842
rect 37924 39976 37976 39982
rect 37924 39918 37976 39924
rect 37936 30802 37964 39918
rect 37924 30796 37976 30802
rect 37924 30738 37976 30744
rect 37924 30660 37976 30666
rect 37924 30602 37976 30608
rect 37936 30394 37964 30602
rect 37924 30388 37976 30394
rect 37924 30330 37976 30336
rect 37924 27872 37976 27878
rect 37924 27814 37976 27820
rect 37936 27538 37964 27814
rect 37924 27532 37976 27538
rect 37924 27474 37976 27480
rect 37660 27118 37872 27146
rect 37660 21554 37688 27118
rect 37740 26920 37792 26926
rect 37740 26862 37792 26868
rect 37648 21548 37700 21554
rect 37648 21490 37700 21496
rect 37648 17196 37700 17202
rect 37648 17138 37700 17144
rect 37556 10668 37608 10674
rect 37556 10610 37608 10616
rect 37464 9580 37516 9586
rect 37464 9522 37516 9528
rect 37660 7410 37688 17138
rect 37648 7404 37700 7410
rect 37648 7346 37700 7352
rect 37752 6914 37780 26862
rect 37924 25696 37976 25702
rect 37924 25638 37976 25644
rect 37936 25362 37964 25638
rect 37924 25356 37976 25362
rect 37924 25298 37976 25304
rect 37832 24608 37884 24614
rect 37832 24550 37884 24556
rect 37844 23254 37872 24550
rect 37924 23520 37976 23526
rect 37924 23462 37976 23468
rect 37832 23248 37884 23254
rect 37832 23190 37884 23196
rect 37936 23186 37964 23462
rect 37924 23180 37976 23186
rect 37924 23122 37976 23128
rect 37832 22432 37884 22438
rect 37832 22374 37884 22380
rect 37844 22098 37872 22374
rect 37832 22092 37884 22098
rect 37832 22034 37884 22040
rect 37832 21480 37884 21486
rect 37832 21422 37884 21428
rect 37844 12918 37872 21422
rect 37924 20256 37976 20262
rect 37924 20198 37976 20204
rect 37936 19922 37964 20198
rect 37924 19916 37976 19922
rect 37924 19858 37976 19864
rect 38028 16114 38056 45766
rect 38106 44296 38162 44305
rect 38106 44231 38162 44240
rect 38120 43858 38148 44231
rect 38108 43852 38160 43858
rect 38108 43794 38160 43800
rect 38108 42628 38160 42634
rect 38108 42570 38160 42576
rect 38120 42265 38148 42570
rect 38106 42256 38162 42265
rect 38106 42191 38162 42200
rect 38212 40594 38240 49286
rect 38630 49200 38742 50000
rect 39274 49200 39386 50000
rect 38384 45484 38436 45490
rect 38384 45426 38436 45432
rect 38396 41002 38424 45426
rect 38384 40996 38436 41002
rect 38384 40938 38436 40944
rect 38200 40588 38252 40594
rect 38200 40530 38252 40536
rect 38200 39840 38252 39846
rect 38200 39782 38252 39788
rect 38106 39536 38162 39545
rect 38106 39471 38108 39480
rect 38160 39471 38162 39480
rect 38108 39442 38160 39448
rect 38212 38418 38240 39782
rect 38200 38412 38252 38418
rect 38200 38354 38252 38360
rect 38106 38176 38162 38185
rect 38106 38111 38162 38120
rect 38120 37330 38148 38111
rect 38292 37868 38344 37874
rect 38292 37810 38344 37816
rect 38108 37324 38160 37330
rect 38108 37266 38160 37272
rect 38108 35624 38160 35630
rect 38108 35566 38160 35572
rect 38120 35465 38148 35566
rect 38106 35456 38162 35465
rect 38106 35391 38162 35400
rect 38108 33856 38160 33862
rect 38108 33798 38160 33804
rect 38120 33590 38148 33798
rect 38108 33584 38160 33590
rect 38108 33526 38160 33532
rect 38106 32056 38162 32065
rect 38106 31991 38162 32000
rect 38120 31890 38148 31991
rect 38108 31884 38160 31890
rect 38108 31826 38160 31832
rect 38200 30728 38252 30734
rect 38200 30670 38252 30676
rect 38106 30016 38162 30025
rect 38106 29951 38162 29960
rect 38120 29714 38148 29951
rect 38108 29708 38160 29714
rect 38108 29650 38160 29656
rect 38212 29170 38240 30670
rect 38200 29164 38252 29170
rect 38200 29106 38252 29112
rect 38108 28552 38160 28558
rect 38108 28494 38160 28500
rect 38120 27538 38148 28494
rect 38108 27532 38160 27538
rect 38108 27474 38160 27480
rect 38108 25696 38160 25702
rect 38108 25638 38160 25644
rect 38120 25362 38148 25638
rect 38108 25356 38160 25362
rect 38108 25298 38160 25304
rect 38106 24576 38162 24585
rect 38106 24511 38162 24520
rect 38120 24274 38148 24511
rect 38108 24268 38160 24274
rect 38108 24210 38160 24216
rect 38304 23730 38332 37810
rect 38396 28150 38424 40938
rect 38476 36780 38528 36786
rect 38476 36722 38528 36728
rect 38384 28144 38436 28150
rect 38384 28086 38436 28092
rect 38292 23724 38344 23730
rect 38292 23666 38344 23672
rect 38488 22094 38516 36722
rect 38212 22066 38516 22094
rect 38106 21176 38162 21185
rect 38106 21111 38162 21120
rect 38120 21010 38148 21111
rect 38108 21004 38160 21010
rect 38108 20946 38160 20952
rect 38212 20466 38240 22066
rect 38200 20460 38252 20466
rect 38200 20402 38252 20408
rect 38108 19848 38160 19854
rect 38108 19790 38160 19796
rect 38120 19378 38148 19790
rect 38108 19372 38160 19378
rect 38108 19314 38160 19320
rect 38108 18692 38160 18698
rect 38108 18634 38160 18640
rect 38120 18465 38148 18634
rect 38106 18456 38162 18465
rect 38106 18391 38162 18400
rect 38106 17776 38162 17785
rect 38106 17711 38108 17720
rect 38160 17711 38162 17720
rect 38108 17682 38160 17688
rect 38106 17096 38162 17105
rect 38106 17031 38162 17040
rect 38120 16658 38148 17031
rect 38108 16652 38160 16658
rect 38108 16594 38160 16600
rect 38016 16108 38068 16114
rect 38016 16050 38068 16056
rect 38106 15736 38162 15745
rect 38106 15671 38162 15680
rect 38120 15570 38148 15671
rect 38108 15564 38160 15570
rect 38108 15506 38160 15512
rect 37832 12912 37884 12918
rect 37832 12854 37884 12860
rect 38108 12844 38160 12850
rect 38108 12786 38160 12792
rect 38120 12345 38148 12786
rect 38106 12336 38162 12345
rect 38106 12271 38162 12280
rect 38108 12232 38160 12238
rect 38108 12174 38160 12180
rect 37924 11552 37976 11558
rect 37924 11494 37976 11500
rect 37936 11218 37964 11494
rect 38120 11218 38148 12174
rect 37924 11212 37976 11218
rect 37924 11154 37976 11160
rect 38108 11212 38160 11218
rect 38108 11154 38160 11160
rect 38108 10464 38160 10470
rect 38108 10406 38160 10412
rect 38016 9988 38068 9994
rect 38016 9930 38068 9936
rect 37924 9376 37976 9382
rect 37924 9318 37976 9324
rect 37936 9042 37964 9318
rect 37924 9036 37976 9042
rect 37924 8978 37976 8984
rect 37832 7880 37884 7886
rect 37832 7822 37884 7828
rect 37384 6886 37504 6914
rect 37372 4616 37424 4622
rect 37372 4558 37424 4564
rect 37280 4140 37332 4146
rect 37280 4082 37332 4088
rect 37280 3936 37332 3942
rect 37280 3878 37332 3884
rect 36636 3188 36688 3194
rect 36636 3130 36688 3136
rect 36648 1578 36676 3130
rect 36728 2372 36780 2378
rect 36728 2314 36780 2320
rect 36740 2145 36768 2314
rect 37292 2310 37320 3878
rect 37384 2582 37412 4558
rect 37476 3602 37504 6886
rect 37660 6886 37780 6914
rect 37556 6316 37608 6322
rect 37556 6258 37608 6264
rect 37464 3596 37516 3602
rect 37464 3538 37516 3544
rect 37464 3460 37516 3466
rect 37464 3402 37516 3408
rect 37476 3194 37504 3402
rect 37464 3188 37516 3194
rect 37464 3130 37516 3136
rect 37568 3126 37596 6258
rect 37556 3120 37608 3126
rect 37556 3062 37608 3068
rect 37660 3058 37688 6886
rect 37844 6338 37872 7822
rect 37924 7200 37976 7206
rect 37924 7142 37976 7148
rect 37936 6866 37964 7142
rect 37924 6860 37976 6866
rect 37924 6802 37976 6808
rect 37752 6310 37872 6338
rect 37752 5846 37780 6310
rect 37832 6248 37884 6254
rect 37832 6190 37884 6196
rect 37740 5840 37792 5846
rect 37740 5782 37792 5788
rect 37844 5234 37872 6190
rect 37924 6112 37976 6118
rect 37924 6054 37976 6060
rect 37936 5778 37964 6054
rect 37924 5772 37976 5778
rect 37924 5714 37976 5720
rect 37832 5228 37884 5234
rect 37832 5170 37884 5176
rect 37648 3052 37700 3058
rect 37648 2994 37700 3000
rect 37372 2576 37424 2582
rect 37372 2518 37424 2524
rect 37280 2304 37332 2310
rect 37280 2246 37332 2252
rect 36726 2136 36782 2145
rect 36726 2071 36782 2080
rect 36648 1550 36768 1578
rect 36740 800 36768 1550
rect 38028 800 38056 9930
rect 38120 9042 38148 10406
rect 38108 9036 38160 9042
rect 38108 8978 38160 8984
rect 38108 8356 38160 8362
rect 38108 8298 38160 8304
rect 38120 6866 38148 8298
rect 38108 6860 38160 6866
rect 38108 6802 38160 6808
rect 38108 3528 38160 3534
rect 38108 3470 38160 3476
rect 38120 2650 38148 3470
rect 38108 2644 38160 2650
rect 38108 2586 38160 2592
rect 35806 776 35862 785
rect 35806 711 35862 720
rect 36054 0 36166 800
rect 36698 0 36810 800
rect 37986 0 38098 800
rect 38630 0 38742 800
rect 39274 0 39386 800
<< via2 >>
rect 2962 49680 3018 49736
rect 1398 47640 1454 47696
rect 1398 44920 1454 44976
rect 1398 41556 1400 41576
rect 1400 41556 1452 41576
rect 1452 41556 1454 41576
rect 1398 41520 1454 41556
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 3330 46960 3386 47016
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 1398 36116 1400 36136
rect 1400 36116 1452 36136
rect 1452 36116 1454 36136
rect 1398 36080 1454 36116
rect 1858 21800 1914 21856
rect 1858 19760 1914 19816
rect 1858 16360 1914 16416
rect 1398 15680 1454 15736
rect 1582 10240 1638 10296
rect 1398 5480 1454 5536
rect 2778 43560 2834 43616
rect 2962 42200 3018 42256
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 2870 38836 2872 38856
rect 2872 38836 2924 38856
rect 2924 38836 2926 38856
rect 2870 38800 2926 38836
rect 2778 29280 2834 29336
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 3422 40840 3478 40896
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 3330 37440 3386 37496
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 2778 22516 2780 22536
rect 2780 22516 2832 22536
rect 2832 22516 2834 22536
rect 2778 22480 2834 22516
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 2778 13640 2834 13696
rect 2778 12960 2834 13016
rect 2778 9560 2834 9616
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 2778 8200 2834 8256
rect 2778 6860 2834 6896
rect 2778 6840 2780 6860
rect 2780 6840 2832 6860
rect 2832 6840 2834 6860
rect 2778 2080 2834 2136
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3974 4800 4030 4856
rect 4066 4120 4122 4176
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 2870 1400 2926 1456
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 6642 3440 6698 3496
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 15658 29572 15714 29608
rect 15658 29552 15660 29572
rect 15660 29552 15712 29572
rect 15712 29552 15714 29572
rect 15658 29044 15660 29064
rect 15660 29044 15712 29064
rect 15712 29044 15714 29064
rect 15658 29008 15714 29044
rect 15934 27956 15936 27976
rect 15936 27956 15988 27976
rect 15988 27956 15990 27976
rect 15934 27920 15990 27956
rect 15842 25916 15844 25936
rect 15844 25916 15896 25936
rect 15896 25916 15898 25936
rect 15842 25880 15898 25916
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 15750 4256 15806 4312
rect 15658 3984 15714 4040
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 23570 35128 23626 35184
rect 25778 35148 25834 35184
rect 25778 35128 25780 35148
rect 25780 35128 25832 35148
rect 25832 35128 25834 35148
rect 35806 49000 35862 49056
rect 35346 47640 35402 47696
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 37094 46280 37150 46336
rect 35806 45600 35862 45656
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 35806 42880 35862 42936
rect 34610 41540 34666 41576
rect 34610 41520 34612 41540
rect 34612 41520 34664 41540
rect 34664 41520 34666 41540
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 37094 40160 37150 40216
rect 37094 38800 37150 38856
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35714 34040 35770 34096
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35806 29280 35862 29336
rect 35346 26560 35402 26616
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 23018 3712 23074 3768
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 37186 30640 37242 30696
rect 37186 27920 37242 27976
rect 37186 25880 37242 25936
rect 37186 23840 37242 23896
rect 37186 21800 37242 21856
rect 37186 20440 37242 20496
rect 37186 11600 37242 11656
rect 37186 9560 37242 9616
rect 37186 7520 37242 7576
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35254 5480 35310 5536
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34610 4120 34666 4176
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35346 2796 35348 2816
rect 35348 2796 35400 2816
rect 35400 2796 35402 2816
rect 35346 2760 35402 2796
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37186 6160 37242 6216
rect 35530 1400 35586 1456
rect 38106 44240 38162 44296
rect 38106 42200 38162 42256
rect 38106 39500 38162 39536
rect 38106 39480 38108 39500
rect 38108 39480 38160 39500
rect 38160 39480 38162 39500
rect 38106 38120 38162 38176
rect 38106 35400 38162 35456
rect 38106 32000 38162 32056
rect 38106 29960 38162 30016
rect 38106 24520 38162 24576
rect 38106 21120 38162 21176
rect 38106 18400 38162 18456
rect 38106 17740 38162 17776
rect 38106 17720 38108 17740
rect 38108 17720 38160 17740
rect 38160 17720 38162 17740
rect 38106 17040 38162 17096
rect 38106 15680 38162 15736
rect 38106 12280 38162 12336
rect 36726 2080 36782 2136
rect 35806 720 35862 776
<< metal3 >>
rect 0 49738 800 49828
rect 2957 49738 3023 49741
rect 0 49736 3023 49738
rect 0 49680 2962 49736
rect 3018 49680 3023 49736
rect 0 49678 3023 49680
rect 0 49588 800 49678
rect 2957 49675 3023 49678
rect 35801 49058 35867 49061
rect 39200 49058 40000 49148
rect 35801 49056 40000 49058
rect 35801 49000 35806 49056
rect 35862 49000 40000 49056
rect 35801 48998 40000 49000
rect 35801 48995 35867 48998
rect 39200 48908 40000 48998
rect 0 48228 800 48468
rect 39200 48228 40000 48468
rect 0 47698 800 47788
rect 1393 47698 1459 47701
rect 0 47696 1459 47698
rect 0 47640 1398 47696
rect 1454 47640 1459 47696
rect 0 47638 1459 47640
rect 0 47548 800 47638
rect 1393 47635 1459 47638
rect 35341 47698 35407 47701
rect 39200 47698 40000 47788
rect 35341 47696 40000 47698
rect 35341 47640 35346 47696
rect 35402 47640 40000 47696
rect 35341 47638 40000 47640
rect 35341 47635 35407 47638
rect 39200 47548 40000 47638
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47108
rect 3325 47018 3391 47021
rect 0 47016 3391 47018
rect 0 46960 3330 47016
rect 3386 46960 3391 47016
rect 0 46958 3391 46960
rect 0 46868 800 46958
rect 3325 46955 3391 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 37089 46338 37155 46341
rect 39200 46338 40000 46428
rect 37089 46336 40000 46338
rect 37089 46280 37094 46336
rect 37150 46280 40000 46336
rect 37089 46278 40000 46280
rect 37089 46275 37155 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 46207 35248 46208
rect 39200 46188 40000 46278
rect 0 45508 800 45748
rect 19568 45728 19888 45729
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 35801 45658 35867 45661
rect 39200 45658 40000 45748
rect 35801 45656 40000 45658
rect 35801 45600 35806 45656
rect 35862 45600 40000 45656
rect 35801 45598 40000 45600
rect 35801 45595 35867 45598
rect 39200 45508 40000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45068
rect 1393 44978 1459 44981
rect 0 44976 1459 44978
rect 0 44920 1398 44976
rect 1454 44920 1459 44976
rect 0 44918 1459 44920
rect 0 44828 800 44918
rect 1393 44915 1459 44918
rect 39200 44828 40000 45068
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 0 44148 800 44388
rect 38101 44298 38167 44301
rect 39200 44298 40000 44388
rect 38101 44296 40000 44298
rect 38101 44240 38106 44296
rect 38162 44240 40000 44296
rect 38101 44238 40000 44240
rect 38101 44235 38167 44238
rect 39200 44148 40000 44238
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43708
rect 2773 43618 2839 43621
rect 0 43616 2839 43618
rect 0 43560 2778 43616
rect 2834 43560 2839 43616
rect 0 43558 2839 43560
rect 0 43468 800 43558
rect 2773 43555 2839 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 43487 19888 43488
rect 4208 43008 4528 43009
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 35801 42938 35867 42941
rect 39200 42938 40000 43028
rect 35801 42936 40000 42938
rect 35801 42880 35806 42936
rect 35862 42880 40000 42936
rect 35801 42878 40000 42880
rect 35801 42875 35867 42878
rect 39200 42788 40000 42878
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 0 42258 800 42348
rect 2957 42258 3023 42261
rect 0 42256 3023 42258
rect 0 42200 2962 42256
rect 3018 42200 3023 42256
rect 0 42198 3023 42200
rect 0 42108 800 42198
rect 2957 42195 3023 42198
rect 38101 42258 38167 42261
rect 39200 42258 40000 42348
rect 38101 42256 40000 42258
rect 38101 42200 38106 42256
rect 38162 42200 40000 42256
rect 38101 42198 40000 42200
rect 38101 42195 38167 42198
rect 39200 42108 40000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41668
rect 1393 41578 1459 41581
rect 0 41576 1459 41578
rect 0 41520 1398 41576
rect 1454 41520 1459 41576
rect 0 41518 1459 41520
rect 0 41428 800 41518
rect 1393 41515 1459 41518
rect 34605 41578 34671 41581
rect 39200 41578 40000 41668
rect 34605 41576 40000 41578
rect 34605 41520 34610 41576
rect 34666 41520 40000 41576
rect 34605 41518 40000 41520
rect 34605 41515 34671 41518
rect 39200 41428 40000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40898 800 40988
rect 3417 40898 3483 40901
rect 0 40896 3483 40898
rect 0 40840 3422 40896
rect 3478 40840 3483 40896
rect 0 40838 3483 40840
rect 0 40748 800 40838
rect 3417 40835 3483 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 40767 35248 40768
rect 0 40068 800 40308
rect 19568 40288 19888 40289
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 37089 40218 37155 40221
rect 39200 40218 40000 40308
rect 37089 40216 40000 40218
rect 37089 40160 37094 40216
rect 37150 40160 40000 40216
rect 37089 40158 40000 40160
rect 37089 40155 37155 40158
rect 39200 40068 40000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 38101 39538 38167 39541
rect 39200 39538 40000 39628
rect 38101 39536 40000 39538
rect 38101 39480 38106 39536
rect 38162 39480 40000 39536
rect 38101 39478 40000 39480
rect 38101 39475 38167 39478
rect 39200 39388 40000 39478
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38858 800 38948
rect 2865 38858 2931 38861
rect 0 38856 2931 38858
rect 0 38800 2870 38856
rect 2926 38800 2931 38856
rect 0 38798 2931 38800
rect 0 38708 800 38798
rect 2865 38795 2931 38798
rect 37089 38858 37155 38861
rect 39200 38858 40000 38948
rect 37089 38856 40000 38858
rect 37089 38800 37094 38856
rect 37150 38800 40000 38856
rect 37089 38798 40000 38800
rect 37089 38795 37155 38798
rect 39200 38708 40000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38028 800 38268
rect 38101 38178 38167 38181
rect 39200 38178 40000 38268
rect 38101 38176 40000 38178
rect 38101 38120 38106 38176
rect 38162 38120 40000 38176
rect 38101 38118 40000 38120
rect 38101 38115 38167 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 38047 19888 38048
rect 39200 38028 40000 38118
rect 0 37498 800 37588
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 3325 37498 3391 37501
rect 0 37496 3391 37498
rect 0 37440 3330 37496
rect 3386 37440 3391 37496
rect 0 37438 3391 37440
rect 0 37348 800 37438
rect 3325 37435 3391 37438
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 39200 36668 40000 36908
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36138 800 36228
rect 1393 36138 1459 36141
rect 0 36136 1459 36138
rect 0 36080 1398 36136
rect 1454 36080 1459 36136
rect 0 36078 1459 36080
rect 0 35988 800 36078
rect 1393 36075 1459 36078
rect 39200 35988 40000 36228
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 0 35308 800 35548
rect 38101 35458 38167 35461
rect 39200 35458 40000 35548
rect 38101 35456 40000 35458
rect 38101 35400 38106 35456
rect 38162 35400 40000 35456
rect 38101 35398 40000 35400
rect 38101 35395 38167 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 35327 35248 35328
rect 39200 35308 40000 35398
rect 23565 35186 23631 35189
rect 25773 35186 25839 35189
rect 23565 35184 25839 35186
rect 23565 35128 23570 35184
rect 23626 35128 25778 35184
rect 25834 35128 25839 35184
rect 23565 35126 25839 35128
rect 23565 35123 23631 35126
rect 25773 35123 25839 35126
rect 0 34628 800 34868
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 33948 800 34188
rect 35709 34098 35775 34101
rect 39200 34098 40000 34188
rect 35709 34096 40000 34098
rect 35709 34040 35714 34096
rect 35770 34040 40000 34096
rect 35709 34038 40000 34040
rect 35709 34035 35775 34038
rect 39200 33948 40000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 39200 33268 40000 33508
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 0 32588 800 32828
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 39200 32588 40000 32828
rect 0 31908 800 32148
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 38101 32058 38167 32061
rect 39200 32058 40000 32148
rect 38101 32056 40000 32058
rect 38101 32000 38106 32056
rect 38162 32000 40000 32056
rect 38101 31998 40000 32000
rect 38101 31995 38167 31998
rect 39200 31908 40000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31228 800 31468
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 37181 30698 37247 30701
rect 39200 30698 40000 30788
rect 37181 30696 40000 30698
rect 37181 30640 37186 30696
rect 37242 30640 40000 30696
rect 37181 30638 40000 30640
rect 37181 30635 37247 30638
rect 39200 30548 40000 30638
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 0 29868 800 30108
rect 38101 30018 38167 30021
rect 39200 30018 40000 30108
rect 38101 30016 40000 30018
rect 38101 29960 38106 30016
rect 38162 29960 40000 30016
rect 38101 29958 40000 29960
rect 38101 29955 38167 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 39200 29868 40000 29958
rect 15510 29548 15516 29612
rect 15580 29610 15586 29612
rect 15653 29610 15719 29613
rect 15580 29608 15719 29610
rect 15580 29552 15658 29608
rect 15714 29552 15719 29608
rect 15580 29550 15719 29552
rect 15580 29548 15586 29550
rect 15653 29547 15719 29550
rect 0 29338 800 29428
rect 19568 29408 19888 29409
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 2773 29338 2839 29341
rect 0 29336 2839 29338
rect 0 29280 2778 29336
rect 2834 29280 2839 29336
rect 0 29278 2839 29280
rect 0 29188 800 29278
rect 2773 29275 2839 29278
rect 35801 29338 35867 29341
rect 39200 29338 40000 29428
rect 35801 29336 40000 29338
rect 35801 29280 35806 29336
rect 35862 29280 40000 29336
rect 35801 29278 40000 29280
rect 35801 29275 35867 29278
rect 39200 29188 40000 29278
rect 15653 29068 15719 29069
rect 15653 29066 15700 29068
rect 15608 29064 15700 29066
rect 15608 29008 15658 29064
rect 15608 29006 15700 29008
rect 15653 29004 15700 29006
rect 15764 29004 15770 29068
rect 15653 29003 15719 29004
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 0 28508 800 28748
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 0 27828 800 28068
rect 15929 27978 15995 27981
rect 16062 27978 16068 27980
rect 15929 27976 16068 27978
rect 15929 27920 15934 27976
rect 15990 27920 16068 27976
rect 15929 27918 16068 27920
rect 15929 27915 15995 27918
rect 16062 27916 16068 27918
rect 16132 27916 16138 27980
rect 37181 27978 37247 27981
rect 39200 27978 40000 28068
rect 37181 27976 40000 27978
rect 37181 27920 37186 27976
rect 37242 27920 40000 27976
rect 37181 27918 40000 27920
rect 37181 27915 37247 27918
rect 39200 27828 40000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 39200 27148 40000 27388
rect 0 26468 800 26708
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 35341 26618 35407 26621
rect 39200 26618 40000 26708
rect 35341 26616 40000 26618
rect 35341 26560 35346 26616
rect 35402 26560 40000 26616
rect 35341 26558 40000 26560
rect 35341 26555 35407 26558
rect 39200 26468 40000 26558
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25788 800 26028
rect 15694 25876 15700 25940
rect 15764 25938 15770 25940
rect 15837 25938 15903 25941
rect 15764 25936 15903 25938
rect 15764 25880 15842 25936
rect 15898 25880 15903 25936
rect 15764 25878 15903 25880
rect 15764 25876 15770 25878
rect 15837 25875 15903 25878
rect 37181 25938 37247 25941
rect 39200 25938 40000 26028
rect 37181 25936 40000 25938
rect 37181 25880 37186 25936
rect 37242 25880 40000 25936
rect 37181 25878 40000 25880
rect 37181 25875 37247 25878
rect 39200 25788 40000 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25108 800 25348
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 38101 24578 38167 24581
rect 39200 24578 40000 24668
rect 38101 24576 40000 24578
rect 38101 24520 38106 24576
rect 38162 24520 40000 24576
rect 38101 24518 40000 24520
rect 38101 24515 38167 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 39200 24428 40000 24518
rect 0 23748 800 23988
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 37181 23898 37247 23901
rect 39200 23898 40000 23988
rect 37181 23896 40000 23898
rect 37181 23840 37186 23896
rect 37242 23840 40000 23896
rect 37181 23838 40000 23840
rect 37181 23835 37247 23838
rect 39200 23748 40000 23838
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23068 800 23308
rect 39200 23068 40000 23308
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22538 800 22628
rect 2773 22538 2839 22541
rect 0 22536 2839 22538
rect 0 22480 2778 22536
rect 2834 22480 2839 22536
rect 0 22478 2839 22480
rect 0 22388 800 22478
rect 2773 22475 2839 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 0 21858 800 21948
rect 1853 21858 1919 21861
rect 0 21856 1919 21858
rect 0 21800 1858 21856
rect 1914 21800 1919 21856
rect 0 21798 1919 21800
rect 0 21708 800 21798
rect 1853 21795 1919 21798
rect 37181 21858 37247 21861
rect 39200 21858 40000 21948
rect 37181 21856 40000 21858
rect 37181 21800 37186 21856
rect 37242 21800 40000 21856
rect 37181 21798 40000 21800
rect 37181 21795 37247 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 39200 21708 40000 21798
rect 4208 21248 4528 21249
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 38101 21178 38167 21181
rect 39200 21178 40000 21268
rect 38101 21176 40000 21178
rect 38101 21120 38106 21176
rect 38162 21120 40000 21176
rect 38101 21118 40000 21120
rect 38101 21115 38167 21118
rect 39200 21028 40000 21118
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20348 800 20588
rect 37181 20498 37247 20501
rect 39200 20498 40000 20588
rect 37181 20496 40000 20498
rect 37181 20440 37186 20496
rect 37242 20440 40000 20496
rect 37181 20438 40000 20440
rect 37181 20435 37247 20438
rect 39200 20348 40000 20438
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 0 19818 800 19908
rect 1853 19818 1919 19821
rect 0 19816 1919 19818
rect 0 19760 1858 19816
rect 1914 19760 1919 19816
rect 0 19758 1919 19760
rect 0 19668 800 19758
rect 1853 19755 1919 19758
rect 39200 19668 40000 19908
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 0 18988 800 19228
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 38101 18458 38167 18461
rect 39200 18458 40000 18548
rect 38101 18456 40000 18458
rect 38101 18400 38106 18456
rect 38162 18400 40000 18456
rect 38101 18398 40000 18400
rect 38101 18395 38167 18398
rect 39200 18308 40000 18398
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 0 17778 800 17868
rect 2773 17778 2839 17781
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 0 17628 800 17718
rect 2773 17715 2839 17718
rect 38101 17778 38167 17781
rect 39200 17778 40000 17868
rect 38101 17776 40000 17778
rect 38101 17720 38106 17776
rect 38162 17720 40000 17776
rect 38101 17718 40000 17720
rect 38101 17715 38167 17718
rect 39200 17628 40000 17718
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 0 16948 800 17188
rect 38101 17098 38167 17101
rect 39200 17098 40000 17188
rect 38101 17096 40000 17098
rect 38101 17040 38106 17096
rect 38162 17040 40000 17096
rect 38101 17038 40000 17040
rect 38101 17035 38167 17038
rect 39200 16948 40000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 0 16418 800 16508
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16268 800 16358
rect 1853 16355 1919 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 0 15738 800 15828
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15588 800 15678
rect 1393 15675 1459 15678
rect 38101 15738 38167 15741
rect 39200 15738 40000 15828
rect 38101 15736 40000 15738
rect 38101 15680 38106 15736
rect 38162 15680 40000 15736
rect 38101 15678 40000 15680
rect 38101 15675 38167 15678
rect 39200 15588 40000 15678
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 39200 14908 40000 15148
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14228 800 14468
rect 39200 14228 40000 14468
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13788
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13548 800 13638
rect 2773 13635 2839 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 39200 13548 40000 13788
rect 0 13018 800 13108
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 2773 13018 2839 13021
rect 0 13016 2839 13018
rect 0 12960 2778 13016
rect 2834 12960 2839 13016
rect 0 12958 2839 12960
rect 0 12868 800 12958
rect 2773 12955 2839 12958
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 38101 12338 38167 12341
rect 39200 12338 40000 12428
rect 38101 12336 40000 12338
rect 38101 12280 38106 12336
rect 38162 12280 40000 12336
rect 38101 12278 40000 12280
rect 38101 12275 38167 12278
rect 39200 12188 40000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11508 800 11748
rect 37181 11658 37247 11661
rect 39200 11658 40000 11748
rect 37181 11656 40000 11658
rect 37181 11600 37186 11656
rect 37242 11600 40000 11656
rect 37181 11598 40000 11600
rect 37181 11595 37247 11598
rect 39200 11508 40000 11598
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 0 10828 800 11068
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 39200 10828 40000 11068
rect 0 10298 800 10388
rect 4208 10368 4528 10369
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 1577 10298 1643 10301
rect 0 10296 1643 10298
rect 0 10240 1582 10296
rect 1638 10240 1643 10296
rect 0 10238 1643 10240
rect 0 10148 800 10238
rect 1577 10235 1643 10238
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9618 800 9708
rect 2773 9618 2839 9621
rect 0 9616 2839 9618
rect 0 9560 2778 9616
rect 2834 9560 2839 9616
rect 0 9558 2839 9560
rect 0 9468 800 9558
rect 2773 9555 2839 9558
rect 37181 9618 37247 9621
rect 39200 9618 40000 9708
rect 37181 9616 40000 9618
rect 37181 9560 37186 9616
rect 37242 9560 40000 9616
rect 37181 9558 40000 9560
rect 37181 9555 37247 9558
rect 39200 9468 40000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 39200 8788 40000 9028
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8258 800 8348
rect 2773 8258 2839 8261
rect 0 8256 2839 8258
rect 0 8200 2778 8256
rect 2834 8200 2839 8256
rect 0 8198 2839 8200
rect 0 8108 800 8198
rect 2773 8195 2839 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 8127 35248 8128
rect 39200 8108 40000 8348
rect 0 7428 800 7668
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 37181 7578 37247 7581
rect 39200 7578 40000 7668
rect 37181 7576 40000 7578
rect 37181 7520 37186 7576
rect 37242 7520 40000 7576
rect 37181 7518 40000 7520
rect 37181 7515 37247 7518
rect 39200 7428 40000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6988
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6748 800 6838
rect 2773 6835 2839 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 37181 6218 37247 6221
rect 39200 6218 40000 6308
rect 37181 6216 40000 6218
rect 37181 6160 37186 6216
rect 37242 6160 40000 6216
rect 37181 6158 40000 6160
rect 37181 6155 37247 6158
rect 39200 6068 40000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5538 800 5628
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5388 800 5478
rect 1393 5475 1459 5478
rect 35249 5538 35315 5541
rect 39200 5538 40000 5628
rect 35249 5536 40000 5538
rect 35249 5480 35254 5536
rect 35310 5480 40000 5536
rect 35249 5478 40000 5480
rect 35249 5475 35315 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 39200 5388 40000 5478
rect 0 4858 800 4948
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 3969 4858 4035 4861
rect 0 4856 4035 4858
rect 0 4800 3974 4856
rect 4030 4800 4035 4856
rect 0 4798 4035 4800
rect 0 4708 800 4798
rect 3969 4795 4035 4798
rect 39200 4708 40000 4948
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 15745 4316 15811 4317
rect 15694 4314 15700 4316
rect 0 4178 800 4268
rect 15654 4254 15700 4314
rect 15764 4312 15811 4316
rect 15806 4256 15811 4312
rect 15694 4252 15700 4254
rect 15764 4252 15811 4256
rect 15745 4251 15811 4252
rect 4061 4178 4127 4181
rect 0 4176 4127 4178
rect 0 4120 4066 4176
rect 4122 4120 4127 4176
rect 0 4118 4127 4120
rect 0 4028 800 4118
rect 4061 4115 4127 4118
rect 34605 4178 34671 4181
rect 39200 4178 40000 4268
rect 34605 4176 40000 4178
rect 34605 4120 34610 4176
rect 34666 4120 40000 4176
rect 34605 4118 40000 4120
rect 34605 4115 34671 4118
rect 15510 3980 15516 4044
rect 15580 4042 15586 4044
rect 15653 4042 15719 4045
rect 15580 4040 15719 4042
rect 15580 3984 15658 4040
rect 15714 3984 15719 4040
rect 39200 4028 40000 4118
rect 15580 3982 15719 3984
rect 15580 3980 15586 3982
rect 15653 3979 15719 3982
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 16062 3708 16068 3772
rect 16132 3770 16138 3772
rect 23013 3770 23079 3773
rect 16132 3768 23079 3770
rect 16132 3712 23018 3768
rect 23074 3712 23079 3768
rect 16132 3710 23079 3712
rect 16132 3708 16138 3710
rect 23013 3707 23079 3710
rect 0 3498 800 3588
rect 6637 3498 6703 3501
rect 0 3496 6703 3498
rect 0 3440 6642 3496
rect 6698 3440 6703 3496
rect 0 3438 6703 3440
rect 0 3348 800 3438
rect 6637 3435 6703 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 35341 2818 35407 2821
rect 39200 2818 40000 2908
rect 35341 2816 40000 2818
rect 35341 2760 35346 2816
rect 35402 2760 40000 2816
rect 35341 2758 40000 2760
rect 35341 2755 35407 2758
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 39200 2668 40000 2758
rect 0 2138 800 2228
rect 19568 2208 19888 2209
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 2773 2138 2839 2141
rect 0 2136 2839 2138
rect 0 2080 2778 2136
rect 2834 2080 2839 2136
rect 0 2078 2839 2080
rect 0 1988 800 2078
rect 2773 2075 2839 2078
rect 36721 2138 36787 2141
rect 39200 2138 40000 2228
rect 36721 2136 40000 2138
rect 36721 2080 36726 2136
rect 36782 2080 40000 2136
rect 36721 2078 40000 2080
rect 36721 2075 36787 2078
rect 39200 1988 40000 2078
rect 0 1458 800 1548
rect 2865 1458 2931 1461
rect 0 1456 2931 1458
rect 0 1400 2870 1456
rect 2926 1400 2931 1456
rect 0 1398 2931 1400
rect 0 1308 800 1398
rect 2865 1395 2931 1398
rect 35525 1458 35591 1461
rect 39200 1458 40000 1548
rect 35525 1456 40000 1458
rect 35525 1400 35530 1456
rect 35586 1400 40000 1456
rect 35525 1398 40000 1400
rect 35525 1395 35591 1398
rect 39200 1308 40000 1398
rect 0 628 800 868
rect 35801 778 35867 781
rect 35801 776 39314 778
rect 35801 720 35806 776
rect 35862 720 39314 776
rect 35801 718 39314 720
rect 35801 715 35867 718
rect 39254 234 39314 718
rect 39070 188 39314 234
rect 39070 174 40000 188
rect 39070 98 39130 174
rect 39200 98 40000 174
rect 39070 38 40000 98
rect 39200 -52 40000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 15516 29548 15580 29612
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 15700 29064 15764 29068
rect 15700 29008 15714 29064
rect 15714 29008 15764 29064
rect 15700 29004 15764 29008
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 16068 27916 16132 27980
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 15700 25876 15764 25940
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 15700 4312 15764 4316
rect 15700 4256 15750 4312
rect 15750 4256 15764 4312
rect 15700 4252 15764 4256
rect 15516 3980 15580 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 16068 3708 16132 3772
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 15515 29612 15581 29613
rect 15515 29548 15516 29612
rect 15580 29548 15581 29612
rect 15515 29547 15581 29548
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 15518 4045 15578 29547
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 15699 29068 15765 29069
rect 15699 29004 15700 29068
rect 15764 29004 15765 29068
rect 15699 29003 15765 29004
rect 15702 25941 15762 29003
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 16067 27980 16133 27981
rect 16067 27916 16068 27980
rect 16132 27916 16133 27980
rect 16067 27915 16133 27916
rect 15699 25940 15765 25941
rect 15699 25876 15700 25940
rect 15764 25876 15765 25940
rect 15699 25875 15765 25876
rect 15702 4317 15762 25875
rect 15699 4316 15765 4317
rect 15699 4252 15700 4316
rect 15764 4252 15765 4316
rect 15699 4251 15765 4252
rect 15515 4044 15581 4045
rect 15515 3980 15516 4044
rect 15580 3980 15581 4044
rect 15515 3979 15581 3980
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 16070 3773 16130 27915
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 16067 3772 16133 3773
rect 16067 3708 16068 3772
rect 16132 3708 16133 3772
rect 16067 3707 16133 3708
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1644511149
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_107
timestamp 1644511149
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1644511149
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1644511149
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1644511149
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_229
timestamp 1644511149
transform 1 0 22172 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_241 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1644511149
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1644511149
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_293
timestamp 1644511149
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1644511149
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_321
timestamp 1644511149
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1644511149
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1644511149
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_400
timestamp 1644511149
transform 1 0 37904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_12
timestamp 1644511149
transform 1 0 2208 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_41
timestamp 1644511149
transform 1 0 4876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_48
timestamp 1644511149
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_81
timestamp 1644511149
transform 1 0 8556 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_106
timestamp 1644511149
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_136
timestamp 1644511149
transform 1 0 13616 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_148
timestamp 1644511149
transform 1 0 14720 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_160
timestamp 1644511149
transform 1 0 15824 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_172
timestamp 1644511149
transform 1 0 16928 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_184
timestamp 1644511149
transform 1 0 18032 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_206
timestamp 1644511149
transform 1 0 20056 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1644511149
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_237
timestamp 1644511149
transform 1 0 22908 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_243
timestamp 1644511149
transform 1 0 23460 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_268
timestamp 1644511149
transform 1 0 25760 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_289
timestamp 1644511149
transform 1 0 27692 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_311
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_323
timestamp 1644511149
transform 1 0 30820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_337
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_370
timestamp 1644511149
transform 1 0 35144 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_378
timestamp 1644511149
transform 1 0 35880 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_382
timestamp 1644511149
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_390
timestamp 1644511149
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_397
timestamp 1644511149
transform 1 0 37628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_3
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_10
timestamp 1644511149
transform 1 0 2024 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_17
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_32
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_59
timestamp 1644511149
transform 1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_66
timestamp 1644511149
transform 1 0 7176 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_74
timestamp 1644511149
transform 1 0 7912 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_79
timestamp 1644511149
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_90
timestamp 1644511149
transform 1 0 9384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_122
timestamp 1644511149
transform 1 0 12328 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_129
timestamp 1644511149
transform 1 0 12972 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 1644511149
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_149
timestamp 1644511149
transform 1 0 14812 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_160
timestamp 1644511149
transform 1 0 15824 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_185
timestamp 1644511149
transform 1 0 18124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_201
timestamp 1644511149
transform 1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_226
timestamp 1644511149
transform 1 0 21896 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_230
timestamp 1644511149
transform 1 0 22264 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1644511149
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1644511149
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_248
timestamp 1644511149
transform 1 0 23920 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_274
timestamp 1644511149
transform 1 0 26312 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_286
timestamp 1644511149
transform 1 0 27416 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_295
timestamp 1644511149
transform 1 0 28244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_302
timestamp 1644511149
transform 1 0 28888 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_333
timestamp 1644511149
transform 1 0 31740 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_341
timestamp 1644511149
transform 1 0 32476 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_346
timestamp 1644511149
transform 1 0 32936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_353
timestamp 1644511149
transform 1 0 33580 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_360
timestamp 1644511149
transform 1 0 34224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_371
timestamp 1644511149
transform 1 0 35236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_378
timestamp 1644511149
transform 1 0 35880 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1644511149
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_30
timestamp 1644511149
transform 1 0 3864 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_38
timestamp 1644511149
transform 1 0 4600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_42
timestamp 1644511149
transform 1 0 4968 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_49
timestamp 1644511149
transform 1 0 5612 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_69
timestamp 1644511149
transform 1 0 7452 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_76
timestamp 1644511149
transform 1 0 8096 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_101
timestamp 1644511149
transform 1 0 10396 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1644511149
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_118
timestamp 1644511149
transform 1 0 11960 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_130
timestamp 1644511149
transform 1 0 13064 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_142
timestamp 1644511149
transform 1 0 14168 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_154
timestamp 1644511149
transform 1 0 15272 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_159
timestamp 1644511149
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1644511149
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_181
timestamp 1644511149
transform 1 0 17756 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_188
timestamp 1644511149
transform 1 0 18400 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_200
timestamp 1644511149
transform 1 0 19504 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_206
timestamp 1644511149
transform 1 0 20056 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_210
timestamp 1644511149
transform 1 0 20424 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_222
timestamp 1644511149
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_232
timestamp 1644511149
transform 1 0 22448 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_240
timestamp 1644511149
transform 1 0 23184 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_263
timestamp 1644511149
transform 1 0 25300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp 1644511149
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_346
timestamp 1644511149
transform 1 0 32936 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_358
timestamp 1644511149
transform 1 0 34040 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1644511149
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_397
timestamp 1644511149
transform 1 0 37628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1644511149
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_8
timestamp 1644511149
transform 1 0 1840 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_23
timestamp 1644511149
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1644511149
transform 1 0 4048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1644511149
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_46
timestamp 1644511149
transform 1 0 5336 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_53
timestamp 1644511149
transform 1 0 5980 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1644511149
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_91
timestamp 1644511149
transform 1 0 9476 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_98
timestamp 1644511149
transform 1 0 10120 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_110
timestamp 1644511149
transform 1 0 11224 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_122
timestamp 1644511149
transform 1 0 12328 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_134
timestamp 1644511149
transform 1 0 13432 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_174
timestamp 1644511149
transform 1 0 17112 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_186
timestamp 1644511149
transform 1 0 18216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1644511149
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_232
timestamp 1644511149
transform 1 0 22448 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_244
timestamp 1644511149
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_321
timestamp 1644511149
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_333
timestamp 1644511149
transform 1 0 31740 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_360
timestamp 1644511149
transform 1 0 34224 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_368
timestamp 1644511149
transform 1 0 34960 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_393
timestamp 1644511149
transform 1 0 37260 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_400
timestamp 1644511149
transform 1 0 37904 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1644511149
transform 1 0 38456 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_11
timestamp 1644511149
transform 1 0 2116 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_19
timestamp 1644511149
transform 1 0 2852 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_41
timestamp 1644511149
transform 1 0 4876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1644511149
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_5_60
timestamp 1644511149
transform 1 0 6624 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_66
timestamp 1644511149
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_70
timestamp 1644511149
transform 1 0 7544 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_82
timestamp 1644511149
transform 1 0 8648 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_94
timestamp 1644511149
transform 1 0 9752 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_106
timestamp 1644511149
transform 1 0 10856 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_346
timestamp 1644511149
transform 1 0 32936 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_350
timestamp 1644511149
transform 1 0 33304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_372
timestamp 1644511149
transform 1 0 35328 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_380
timestamp 1644511149
transform 1 0 36064 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_384
timestamp 1644511149
transform 1 0 36432 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_396
timestamp 1644511149
transform 1 0 37536 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1644511149
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1644511149
transform 1 0 3312 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_265
timestamp 1644511149
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_277
timestamp 1644511149
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_289
timestamp 1644511149
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1644511149
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_354
timestamp 1644511149
transform 1 0 33672 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1644511149
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_370
timestamp 1644511149
transform 1 0 35144 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_381
timestamp 1644511149
transform 1 0 36156 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1644511149
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_12
timestamp 1644511149
transform 1 0 2208 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_19
timestamp 1644511149
transform 1 0 2852 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_31
timestamp 1644511149
transform 1 0 3956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_43
timestamp 1644511149
transform 1 0 5060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1644511149
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_249
timestamp 1644511149
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_261
timestamp 1644511149
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1644511149
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_388
timestamp 1644511149
transform 1 0 36800 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_398
timestamp 1644511149
transform 1 0 37720 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_406
timestamp 1644511149
transform 1 0 38456 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_265
timestamp 1644511149
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_277
timestamp 1644511149
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_333
timestamp 1644511149
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_345
timestamp 1644511149
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1644511149
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1644511149
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_381
timestamp 1644511149
transform 1 0 36156 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1644511149
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_14
timestamp 1644511149
transform 1 0 2392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_26
timestamp 1644511149
transform 1 0 3496 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_38
timestamp 1644511149
transform 1 0 4600 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_50
timestamp 1644511149
transform 1 0 5704 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_193
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_205
timestamp 1644511149
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1644511149
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1644511149
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_237
timestamp 1644511149
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_249
timestamp 1644511149
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1644511149
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_305
timestamp 1644511149
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_317
timestamp 1644511149
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1644511149
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_398
timestamp 1644511149
transform 1 0 37720 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_406
timestamp 1644511149
transform 1 0 38456 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1644511149
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_209
timestamp 1644511149
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_221
timestamp 1644511149
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_233
timestamp 1644511149
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1644511149
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1644511149
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_289
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1644511149
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1644511149
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_321
timestamp 1644511149
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_333
timestamp 1644511149
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_345
timestamp 1644511149
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1644511149
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_10_400
timestamp 1644511149
transform 1 0 37904 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1644511149
transform 1 0 38456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_6
timestamp 1644511149
transform 1 0 1656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_31
timestamp 1644511149
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_43
timestamp 1644511149
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_193
timestamp 1644511149
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_205
timestamp 1644511149
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1644511149
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1644511149
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_305
timestamp 1644511149
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_317
timestamp 1644511149
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_400
timestamp 1644511149
transform 1 0 37904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_406
timestamp 1644511149
transform 1 0 38456 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_7
timestamp 1644511149
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_11
timestamp 1644511149
transform 1 0 2116 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_18
timestamp 1644511149
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1644511149
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_177
timestamp 1644511149
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1644511149
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1644511149
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_209
timestamp 1644511149
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_221
timestamp 1644511149
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_233
timestamp 1644511149
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1644511149
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_277
timestamp 1644511149
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_289
timestamp 1644511149
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1644511149
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_381
timestamp 1644511149
transform 1 0 36156 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1644511149
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_7
timestamp 1644511149
transform 1 0 1748 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_29
timestamp 1644511149
transform 1 0 3772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_41
timestamp 1644511149
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1644511149
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_193
timestamp 1644511149
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_205
timestamp 1644511149
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1644511149
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_249
timestamp 1644511149
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_261
timestamp 1644511149
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1644511149
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1644511149
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1644511149
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_305
timestamp 1644511149
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_317
timestamp 1644511149
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1644511149
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_388
timestamp 1644511149
transform 1 0 36800 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_398
timestamp 1644511149
transform 1 0 37720 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_406
timestamp 1644511149
transform 1 0 38456 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_9
timestamp 1644511149
transform 1 0 1932 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_16
timestamp 1644511149
transform 1 0 2576 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_197
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_209
timestamp 1644511149
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_221
timestamp 1644511149
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_233
timestamp 1644511149
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1644511149
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1644511149
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_265
timestamp 1644511149
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1644511149
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_321
timestamp 1644511149
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_333
timestamp 1644511149
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_345
timestamp 1644511149
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1644511149
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_381
timestamp 1644511149
transform 1 0 36156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_403
timestamp 1644511149
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_26
timestamp 1644511149
transform 1 0 3496 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_38
timestamp 1644511149
transform 1 0 4600 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_50
timestamp 1644511149
transform 1 0 5704 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_205
timestamp 1644511149
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1644511149
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_249
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_261
timestamp 1644511149
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1644511149
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1644511149
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1644511149
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_305
timestamp 1644511149
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_317
timestamp 1644511149
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1644511149
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1644511149
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_396
timestamp 1644511149
transform 1 0 37536 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1644511149
transform 1 0 38180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_7
timestamp 1644511149
transform 1 0 1748 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_11
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_18
timestamp 1644511149
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1644511149
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_177
timestamp 1644511149
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1644511149
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_233
timestamp 1644511149
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1644511149
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_265
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_277
timestamp 1644511149
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_289
timestamp 1644511149
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1644511149
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_321
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1644511149
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1644511149
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_381
timestamp 1644511149
transform 1 0 36156 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1644511149
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1644511149
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1644511149
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1644511149
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1644511149
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_181
timestamp 1644511149
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_193
timestamp 1644511149
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_205
timestamp 1644511149
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1644511149
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_237
timestamp 1644511149
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_249
timestamp 1644511149
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_261
timestamp 1644511149
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1644511149
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_305
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_317
timestamp 1644511149
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1644511149
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1644511149
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_397
timestamp 1644511149
transform 1 0 37628 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1644511149
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_13
timestamp 1644511149
transform 1 0 2300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1644511149
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1644511149
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1644511149
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_209
timestamp 1644511149
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_221
timestamp 1644511149
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_233
timestamp 1644511149
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1644511149
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_265
timestamp 1644511149
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_277
timestamp 1644511149
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_289
timestamp 1644511149
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1644511149
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1644511149
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_309
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_321
timestamp 1644511149
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_333
timestamp 1644511149
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_345
timestamp 1644511149
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1644511149
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1644511149
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_18_400
timestamp 1644511149
transform 1 0 37904 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1644511149
transform 1 0 38456 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_3
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1644511149
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1644511149
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1644511149
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_181
timestamp 1644511149
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_193
timestamp 1644511149
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_205
timestamp 1644511149
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1644511149
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_237
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_249
timestamp 1644511149
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1644511149
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1644511149
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1644511149
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_305
timestamp 1644511149
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1644511149
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_403
timestamp 1644511149
transform 1 0 38180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_6
timestamp 1644511149
transform 1 0 1656 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_13
timestamp 1644511149
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1644511149
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1644511149
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1644511149
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_197
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_209
timestamp 1644511149
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_221
timestamp 1644511149
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_233
timestamp 1644511149
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_265
timestamp 1644511149
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_277
timestamp 1644511149
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1644511149
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1644511149
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_321
timestamp 1644511149
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_333
timestamp 1644511149
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_345
timestamp 1644511149
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1644511149
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1644511149
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1644511149
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1644511149
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1644511149
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_181
timestamp 1644511149
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_193
timestamp 1644511149
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_205
timestamp 1644511149
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1644511149
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_261
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1644511149
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1644511149
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1644511149
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_305
timestamp 1644511149
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_317
timestamp 1644511149
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1644511149
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1644511149
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_349
timestamp 1644511149
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_361
timestamp 1644511149
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_373
timestamp 1644511149
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1644511149
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1644511149
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_10
timestamp 1644511149
transform 1 0 2024 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_22
timestamp 1644511149
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_209
timestamp 1644511149
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1644511149
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_265
timestamp 1644511149
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_277
timestamp 1644511149
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_289
timestamp 1644511149
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1644511149
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_321
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_333
timestamp 1644511149
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_345
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1644511149
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1644511149
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_11
timestamp 1644511149
transform 1 0 2116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_23
timestamp 1644511149
transform 1 0 3220 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_35
timestamp 1644511149
transform 1 0 4324 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_47
timestamp 1644511149
transform 1 0 5428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1644511149
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_205
timestamp 1644511149
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1644511149
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_249
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1644511149
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1644511149
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_317
timestamp 1644511149
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1644511149
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_349
timestamp 1644511149
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_361
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_373
timestamp 1644511149
transform 1 0 35420 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_381
timestamp 1644511149
transform 1 0 36156 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_387
timestamp 1644511149
transform 1 0 36708 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1644511149
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_24
timestamp 1644511149
transform 1 0 3312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_109
timestamp 1644511149
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_121
timestamp 1644511149
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1644511149
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1644511149
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_177
timestamp 1644511149
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1644511149
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1644511149
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_209
timestamp 1644511149
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_221
timestamp 1644511149
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1644511149
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_265
timestamp 1644511149
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_321
timestamp 1644511149
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_345
timestamp 1644511149
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1644511149
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1644511149
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_381
timestamp 1644511149
transform 1 0 36156 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_403
timestamp 1644511149
transform 1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_12
timestamp 1644511149
transform 1 0 2208 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_19
timestamp 1644511149
transform 1 0 2852 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_31
timestamp 1644511149
transform 1 0 3956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_43
timestamp 1644511149
transform 1 0 5060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_149
timestamp 1644511149
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1644511149
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1644511149
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_181
timestamp 1644511149
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_205
timestamp 1644511149
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1644511149
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1644511149
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_237
timestamp 1644511149
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_249
timestamp 1644511149
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_261
timestamp 1644511149
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1644511149
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_305
timestamp 1644511149
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_317
timestamp 1644511149
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1644511149
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1644511149
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_349
timestamp 1644511149
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_361
timestamp 1644511149
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_373
timestamp 1644511149
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_388
timestamp 1644511149
transform 1 0 36800 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_398
timestamp 1644511149
transform 1 0 37720 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_406
timestamp 1644511149
transform 1 0 38456 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_41
timestamp 1644511149
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_53
timestamp 1644511149
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_65
timestamp 1644511149
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1644511149
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_109
timestamp 1644511149
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_121
timestamp 1644511149
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1644511149
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_165
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_177
timestamp 1644511149
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1644511149
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1644511149
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_221
timestamp 1644511149
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_233
timestamp 1644511149
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1644511149
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1644511149
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_277
timestamp 1644511149
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_289
timestamp 1644511149
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1644511149
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1644511149
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_321
timestamp 1644511149
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_333
timestamp 1644511149
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_345
timestamp 1644511149
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1644511149
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1644511149
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_381
timestamp 1644511149
transform 1 0 36156 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_403
timestamp 1644511149
transform 1 0 38180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_6
timestamp 1644511149
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_13
timestamp 1644511149
transform 1 0 2300 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_25
timestamp 1644511149
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_37
timestamp 1644511149
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1644511149
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_93
timestamp 1644511149
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1644511149
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1644511149
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_149
timestamp 1644511149
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1644511149
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_193
timestamp 1644511149
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_205
timestamp 1644511149
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1644511149
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1644511149
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_249
timestamp 1644511149
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_261
timestamp 1644511149
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_305
timestamp 1644511149
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_317
timestamp 1644511149
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1644511149
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_349
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_361
timestamp 1644511149
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_373
timestamp 1644511149
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1644511149
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_398
timestamp 1644511149
transform 1 0 37720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_406
timestamp 1644511149
transform 1 0 38456 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1644511149
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1644511149
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_85
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1644511149
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_109
timestamp 1644511149
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_121
timestamp 1644511149
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1644511149
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1644511149
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_153
timestamp 1644511149
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_165
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_177
timestamp 1644511149
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_209
timestamp 1644511149
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_233
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1644511149
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1644511149
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_265
timestamp 1644511149
transform 1 0 25484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_284
timestamp 1644511149
transform 1 0 27232 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_296
timestamp 1644511149
transform 1 0 28336 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_315
timestamp 1644511149
transform 1 0 30084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_332
timestamp 1644511149
transform 1 0 31648 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_344
timestamp 1644511149
transform 1 0 32752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_351
timestamp 1644511149
transform 1 0 33396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_381
timestamp 1644511149
transform 1 0 36156 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_403
timestamp 1644511149
transform 1 0 38180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_9
timestamp 1644511149
transform 1 0 1932 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_21
timestamp 1644511149
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_33
timestamp 1644511149
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1644511149
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1644511149
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_81
timestamp 1644511149
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_93
timestamp 1644511149
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1644511149
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1644511149
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_125
timestamp 1644511149
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_137
timestamp 1644511149
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_149
timestamp 1644511149
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1644511149
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_189
timestamp 1644511149
transform 1 0 18492 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_197
timestamp 1644511149
transform 1 0 19228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_202
timestamp 1644511149
transform 1 0 19688 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_214
timestamp 1644511149
transform 1 0 20792 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1644511149
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_237
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_249
timestamp 1644511149
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_261
timestamp 1644511149
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1644511149
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_293
timestamp 1644511149
transform 1 0 28060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_313
timestamp 1644511149
transform 1 0 29900 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_325
timestamp 1644511149
transform 1 0 31004 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_345
timestamp 1644511149
transform 1 0 32844 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_362
timestamp 1644511149
transform 1 0 34408 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_374
timestamp 1644511149
transform 1 0 35512 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_381
timestamp 1644511149
transform 1 0 36156 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_388
timestamp 1644511149
transform 1 0 36800 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_398
timestamp 1644511149
transform 1 0 37720 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_406
timestamp 1644511149
transform 1 0 38456 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_65
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1644511149
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_109
timestamp 1644511149
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_121
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_177
timestamp 1644511149
transform 1 0 17388 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_184
timestamp 1644511149
transform 1 0 18032 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_191
timestamp 1644511149
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_200
timestamp 1644511149
transform 1 0 19504 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_216
timestamp 1644511149
transform 1 0 20976 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_234
timestamp 1644511149
transform 1 0 22632 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_242
timestamp 1644511149
transform 1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1644511149
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_265
timestamp 1644511149
transform 1 0 25484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_273
timestamp 1644511149
transform 1 0 26220 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_281
timestamp 1644511149
transform 1 0 26956 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_294
timestamp 1644511149
transform 1 0 28152 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_313
timestamp 1644511149
transform 1 0 29900 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_321
timestamp 1644511149
transform 1 0 30636 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_326
timestamp 1644511149
transform 1 0 31096 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_337
timestamp 1644511149
transform 1 0 32108 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_348
timestamp 1644511149
transform 1 0 33120 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1644511149
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_372
timestamp 1644511149
transform 1 0 35328 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_380
timestamp 1644511149
transform 1 0 36064 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1644511149
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_11
timestamp 1644511149
transform 1 0 2116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_23
timestamp 1644511149
transform 1 0 3220 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_35
timestamp 1644511149
transform 1 0 4324 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_47
timestamp 1644511149
transform 1 0 5428 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_81
timestamp 1644511149
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1644511149
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1644511149
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_125
timestamp 1644511149
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_137
timestamp 1644511149
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_149
timestamp 1644511149
transform 1 0 14812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_153
timestamp 1644511149
transform 1 0 15180 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_160
timestamp 1644511149
transform 1 0 15824 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1644511149
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_200
timestamp 1644511149
transform 1 0 19504 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_241
timestamp 1644511149
transform 1 0 23276 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_261
timestamp 1644511149
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_276
timestamp 1644511149
transform 1 0 26496 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_286
timestamp 1644511149
transform 1 0 27416 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_308
timestamp 1644511149
transform 1 0 29440 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_320
timestamp 1644511149
transform 1 0 30544 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_349
timestamp 1644511149
transform 1 0 33212 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_357
timestamp 1644511149
transform 1 0 33948 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_365
timestamp 1644511149
transform 1 0 34684 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_377
timestamp 1644511149
transform 1 0 35788 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_389
timestamp 1644511149
transform 1 0 36892 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_400
timestamp 1644511149
transform 1 0 37904 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1644511149
transform 1 0 38456 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1644511149
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1644511149
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_109
timestamp 1644511149
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_121
timestamp 1644511149
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1644511149
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1644511149
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_141
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_158
timestamp 1644511149
transform 1 0 15640 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_178
timestamp 1644511149
transform 1 0 17480 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_187
timestamp 1644511149
transform 1 0 18308 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1644511149
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_205
timestamp 1644511149
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_213
timestamp 1644511149
transform 1 0 20700 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_229
timestamp 1644511149
transform 1 0 22172 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_243
timestamp 1644511149
transform 1 0 23460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_261
timestamp 1644511149
transform 1 0 25116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_273
timestamp 1644511149
transform 1 0 26220 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_296
timestamp 1644511149
transform 1 0 28336 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_313
timestamp 1644511149
transform 1 0 29900 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_324
timestamp 1644511149
transform 1 0 30912 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_336
timestamp 1644511149
transform 1 0 32016 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_341
timestamp 1644511149
transform 1 0 32476 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_353
timestamp 1644511149
transform 1 0 33580 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_361
timestamp 1644511149
transform 1 0 34316 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_365
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_381
timestamp 1644511149
transform 1 0 36156 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1644511149
transform 1 0 38180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_8
timestamp 1644511149
transform 1 0 1840 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_20
timestamp 1644511149
transform 1 0 2944 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_32
timestamp 1644511149
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_44
timestamp 1644511149
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_73
timestamp 1644511149
transform 1 0 7820 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_94
timestamp 1644511149
transform 1 0 9752 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_106
timestamp 1644511149
transform 1 0 10856 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_137
timestamp 1644511149
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1644511149
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_172
timestamp 1644511149
transform 1 0 16928 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_182
timestamp 1644511149
transform 1 0 17848 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_194
timestamp 1644511149
transform 1 0 18952 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_206
timestamp 1644511149
transform 1 0 20056 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_218
timestamp 1644511149
transform 1 0 21160 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_233
timestamp 1644511149
transform 1 0 22540 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_240
timestamp 1644511149
transform 1 0 23184 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_248
timestamp 1644511149
transform 1 0 23920 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_276
timestamp 1644511149
transform 1 0 26496 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_284
timestamp 1644511149
transform 1 0 27232 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_296
timestamp 1644511149
transform 1 0 28336 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_302
timestamp 1644511149
transform 1 0 28888 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_308
timestamp 1644511149
transform 1 0 29440 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1644511149
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_321
timestamp 1644511149
transform 1 0 30636 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1644511149
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1644511149
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_348
timestamp 1644511149
transform 1 0 33120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_356
timestamp 1644511149
transform 1 0 33856 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_366
timestamp 1644511149
transform 1 0 34776 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_378
timestamp 1644511149
transform 1 0 35880 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_384
timestamp 1644511149
transform 1 0 36432 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_388
timestamp 1644511149
transform 1 0 36800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_397
timestamp 1644511149
transform 1 0 37628 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_9
timestamp 1644511149
transform 1 0 1932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_21
timestamp 1644511149
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_65
timestamp 1644511149
transform 1 0 7084 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_73
timestamp 1644511149
transform 1 0 7820 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_80
timestamp 1644511149
transform 1 0 8464 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_93
timestamp 1644511149
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_97
timestamp 1644511149
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_109
timestamp 1644511149
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_121
timestamp 1644511149
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_153
timestamp 1644511149
transform 1 0 15180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_161
timestamp 1644511149
transform 1 0 15916 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_170
timestamp 1644511149
transform 1 0 16744 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_182
timestamp 1644511149
transform 1 0 17848 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1644511149
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_210
timestamp 1644511149
transform 1 0 20424 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_222
timestamp 1644511149
transform 1 0 21528 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1644511149
transform 1 0 22632 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1644511149
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_253
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_265
timestamp 1644511149
transform 1 0 25484 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_273
timestamp 1644511149
transform 1 0 26220 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_279
timestamp 1644511149
transform 1 0 26772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1644511149
transform 1 0 27600 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_299
timestamp 1644511149
transform 1 0 28612 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_322
timestamp 1644511149
transform 1 0 30728 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_335
timestamp 1644511149
transform 1 0 31924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1644511149
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_373
timestamp 1644511149
transform 1 0 35420 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_381
timestamp 1644511149
transform 1 0 36156 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_403
timestamp 1644511149
transform 1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_12
timestamp 1644511149
transform 1 0 2208 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_24
timestamp 1644511149
transform 1 0 3312 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_36
timestamp 1644511149
transform 1 0 4416 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_48
timestamp 1644511149
transform 1 0 5520 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_69
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_73
timestamp 1644511149
transform 1 0 7820 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1644511149
transform 1 0 9016 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_98
timestamp 1644511149
transform 1 0 10120 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1644511149
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_113
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_125
timestamp 1644511149
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_137
timestamp 1644511149
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_149
timestamp 1644511149
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_181
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_196
timestamp 1644511149
transform 1 0 19136 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_207
timestamp 1644511149
transform 1 0 20148 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_211
timestamp 1644511149
transform 1 0 20516 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1644511149
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_234
timestamp 1644511149
transform 1 0 22632 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_238
timestamp 1644511149
transform 1 0 23000 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_255
timestamp 1644511149
transform 1 0 24564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_259
timestamp 1644511149
transform 1 0 24932 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_276
timestamp 1644511149
transform 1 0 26496 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_286
timestamp 1644511149
transform 1 0 27416 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_293
timestamp 1644511149
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_301
timestamp 1644511149
transform 1 0 28796 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_309
timestamp 1644511149
transform 1 0 29532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_313
timestamp 1644511149
transform 1 0 29900 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_324
timestamp 1644511149
transform 1 0 30912 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_344
timestamp 1644511149
transform 1 0 32752 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_351
timestamp 1644511149
transform 1 0 33396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_359
timestamp 1644511149
transform 1 0 34132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_365
timestamp 1644511149
transform 1 0 34684 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1644511149
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_397
timestamp 1644511149
transform 1 0 37628 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1644511149
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1644511149
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_109
timestamp 1644511149
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_121
timestamp 1644511149
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1644511149
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_153
timestamp 1644511149
transform 1 0 15180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_157
timestamp 1644511149
transform 1 0 15548 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_179
timestamp 1644511149
transform 1 0 17572 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_191
timestamp 1644511149
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1644511149
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_205
timestamp 1644511149
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_214
timestamp 1644511149
transform 1 0 20792 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_226
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_236
timestamp 1644511149
transform 1 0 22816 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_243
timestamp 1644511149
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1644511149
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_253
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_273
timestamp 1644511149
transform 1 0 26220 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_280
timestamp 1644511149
transform 1 0 26864 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_292
timestamp 1644511149
transform 1 0 27968 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_297
timestamp 1644511149
transform 1 0 28428 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_305
timestamp 1644511149
transform 1 0 29164 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_321
timestamp 1644511149
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_333
timestamp 1644511149
transform 1 0 31740 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_340
timestamp 1644511149
transform 1 0 32384 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_352
timestamp 1644511149
transform 1 0 33488 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_365
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_378
timestamp 1644511149
transform 1 0 35880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1644511149
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_28
timestamp 1644511149
transform 1 0 3680 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_40
timestamp 1644511149
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_52
timestamp 1644511149
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_149
timestamp 1644511149
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1644511149
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_172
timestamp 1644511149
transform 1 0 16928 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_180
timestamp 1644511149
transform 1 0 17664 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_198
timestamp 1644511149
transform 1 0 19320 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1644511149
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1644511149
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_225
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_233
timestamp 1644511149
transform 1 0 22540 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_240
timestamp 1644511149
transform 1 0 23184 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_247
timestamp 1644511149
transform 1 0 23828 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_258
timestamp 1644511149
transform 1 0 24840 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_270
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1644511149
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_293
timestamp 1644511149
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_304
timestamp 1644511149
transform 1 0 29072 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_317
timestamp 1644511149
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1644511149
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_345
timestamp 1644511149
transform 1 0 32844 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_353
timestamp 1644511149
transform 1 0 33580 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_364
timestamp 1644511149
transform 1 0 34592 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_376
timestamp 1644511149
transform 1 0 35696 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_384
timestamp 1644511149
transform 1 0 36432 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_400
timestamp 1644511149
transform 1 0 37904 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_406
timestamp 1644511149
transform 1 0 38456 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_8
timestamp 1644511149
transform 1 0 1840 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1644511149
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1644511149
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_97
timestamp 1644511149
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_109
timestamp 1644511149
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_121
timestamp 1644511149
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1644511149
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1644511149
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_161
timestamp 1644511149
transform 1 0 15916 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_168
timestamp 1644511149
transform 1 0 16560 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_180
timestamp 1644511149
transform 1 0 17664 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1644511149
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_200
timestamp 1644511149
transform 1 0 19504 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_212
timestamp 1644511149
transform 1 0 20608 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_220
timestamp 1644511149
transform 1 0 21344 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_224
timestamp 1644511149
transform 1 0 21712 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_231
timestamp 1644511149
transform 1 0 22356 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_243
timestamp 1644511149
transform 1 0 23460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1644511149
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_269
timestamp 1644511149
transform 1 0 25852 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_281
timestamp 1644511149
transform 1 0 26956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_287
timestamp 1644511149
transform 1 0 27508 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_295
timestamp 1644511149
transform 1 0 28244 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_318
timestamp 1644511149
transform 1 0 30360 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_326
timestamp 1644511149
transform 1 0 31096 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_343
timestamp 1644511149
transform 1 0 32660 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_351
timestamp 1644511149
transform 1 0 33396 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_356
timestamp 1644511149
transform 1 0 33856 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_375
timestamp 1644511149
transform 1 0 35604 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_381
timestamp 1644511149
transform 1 0 36156 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1644511149
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1644511149
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1644511149
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1644511149
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_69
timestamp 1644511149
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_93
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_125
timestamp 1644511149
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_137
timestamp 1644511149
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_155
timestamp 1644511149
transform 1 0 15364 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_163
timestamp 1644511149
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_169
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_173
timestamp 1644511149
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_200
timestamp 1644511149
transform 1 0 19504 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_212
timestamp 1644511149
transform 1 0 20608 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_218
timestamp 1644511149
transform 1 0 21160 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_39_247
timestamp 1644511149
transform 1 0 23828 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_259
timestamp 1644511149
transform 1 0 24932 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_284
timestamp 1644511149
transform 1 0 27232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_294
timestamp 1644511149
transform 1 0 28152 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_301
timestamp 1644511149
transform 1 0 28796 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_307
timestamp 1644511149
transform 1 0 29348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_317
timestamp 1644511149
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_345
timestamp 1644511149
transform 1 0 32844 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_355
timestamp 1644511149
transform 1 0 33764 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_362
timestamp 1644511149
transform 1 0 34408 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_370
timestamp 1644511149
transform 1 0 35144 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_387
timestamp 1644511149
transform 1 0 36708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1644511149
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_397
timestamp 1644511149
transform 1 0 37628 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_97
timestamp 1644511149
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_109
timestamp 1644511149
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_121
timestamp 1644511149
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1644511149
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_161
timestamp 1644511149
transform 1 0 15916 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_170
timestamp 1644511149
transform 1 0 16744 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_182
timestamp 1644511149
transform 1 0 17848 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1644511149
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_205
timestamp 1644511149
transform 1 0 19964 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_211
timestamp 1644511149
transform 1 0 20516 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_221
timestamp 1644511149
transform 1 0 21436 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_225
timestamp 1644511149
transform 1 0 21804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_235
timestamp 1644511149
transform 1 0 22724 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_247
timestamp 1644511149
transform 1 0 23828 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_265
timestamp 1644511149
transform 1 0 25484 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_40_271
timestamp 1644511149
transform 1 0 26036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_281
timestamp 1644511149
transform 1 0 26956 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1644511149
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1644511149
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_317
timestamp 1644511149
transform 1 0 30268 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_325
timestamp 1644511149
transform 1 0 31004 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_337
timestamp 1644511149
transform 1 0 32108 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_349
timestamp 1644511149
transform 1 0 33212 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_360
timestamp 1644511149
transform 1 0 34224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_365
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_377
timestamp 1644511149
transform 1 0 35788 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_381
timestamp 1644511149
transform 1 0 36156 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1644511149
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_81
timestamp 1644511149
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_93
timestamp 1644511149
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1644511149
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_149
timestamp 1644511149
transform 1 0 14812 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_157
timestamp 1644511149
transform 1 0 15548 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1644511149
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_201
timestamp 1644511149
transform 1 0 19596 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_206
timestamp 1644511149
transform 1 0 20056 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1644511149
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_230
timestamp 1644511149
transform 1 0 22264 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_242
timestamp 1644511149
transform 1 0 23368 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_250
timestamp 1644511149
transform 1 0 24104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_256
timestamp 1644511149
transform 1 0 24656 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_268
timestamp 1644511149
transform 1 0 25760 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_289
timestamp 1644511149
transform 1 0 27692 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_294
timestamp 1644511149
transform 1 0 28152 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_301
timestamp 1644511149
transform 1 0 28796 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_313
timestamp 1644511149
transform 1 0 29900 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_325
timestamp 1644511149
transform 1 0 31004 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_333
timestamp 1644511149
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_340
timestamp 1644511149
transform 1 0 32384 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_346
timestamp 1644511149
transform 1 0 32936 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_350
timestamp 1644511149
transform 1 0 33304 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_360
timestamp 1644511149
transform 1 0 34224 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_369
timestamp 1644511149
transform 1 0 35052 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_373
timestamp 1644511149
transform 1 0 35420 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_381
timestamp 1644511149
transform 1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1644511149
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_400
timestamp 1644511149
transform 1 0 37904 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_406
timestamp 1644511149
transform 1 0 38456 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1644511149
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1644511149
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_97
timestamp 1644511149
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_109
timestamp 1644511149
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_121
timestamp 1644511149
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1644511149
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1644511149
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_153
timestamp 1644511149
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_165
timestamp 1644511149
transform 1 0 16284 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_171
timestamp 1644511149
transform 1 0 16836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_183
timestamp 1644511149
transform 1 0 17940 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 1644511149
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_200
timestamp 1644511149
transform 1 0 19504 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_208
timestamp 1644511149
transform 1 0 20240 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_218
timestamp 1644511149
transform 1 0 21160 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_230
timestamp 1644511149
transform 1 0 22264 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_242
timestamp 1644511149
transform 1 0 23368 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1644511149
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_269
timestamp 1644511149
transform 1 0 25852 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_281
timestamp 1644511149
transform 1 0 26956 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_293
timestamp 1644511149
transform 1 0 28060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1644511149
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_321
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_339
timestamp 1644511149
transform 1 0 32292 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_351
timestamp 1644511149
transform 1 0 33396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_372
timestamp 1644511149
transform 1 0 35328 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_380
timestamp 1644511149
transform 1 0 36064 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_403
timestamp 1644511149
transform 1 0 38180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_69
timestamp 1644511149
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_81
timestamp 1644511149
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_93
timestamp 1644511149
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1644511149
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_113
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_125
timestamp 1644511149
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_137
timestamp 1644511149
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_149
timestamp 1644511149
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1644511149
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_174
timestamp 1644511149
transform 1 0 17112 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_182
timestamp 1644511149
transform 1 0 17848 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_191
timestamp 1644511149
transform 1 0 18676 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_201
timestamp 1644511149
transform 1 0 19596 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_216
timestamp 1644511149
transform 1 0 20976 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_43_228
timestamp 1644511149
transform 1 0 22080 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_234
timestamp 1644511149
transform 1 0 22632 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_241
timestamp 1644511149
transform 1 0 23276 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_253
timestamp 1644511149
transform 1 0 24380 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_259
timestamp 1644511149
transform 1 0 24932 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_270
timestamp 1644511149
transform 1 0 25944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1644511149
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1644511149
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_321
timestamp 1644511149
transform 1 0 30636 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_331
timestamp 1644511149
transform 1 0 31556 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_344
timestamp 1644511149
transform 1 0 32752 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_351
timestamp 1644511149
transform 1 0 33396 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_359
timestamp 1644511149
transform 1 0 34132 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_366
timestamp 1644511149
transform 1 0 34776 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_388
timestamp 1644511149
transform 1 0 36800 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_396
timestamp 1644511149
transform 1 0 37536 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1644511149
transform 1 0 38180 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1644511149
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_65
timestamp 1644511149
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1644511149
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1644511149
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_109
timestamp 1644511149
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_121
timestamp 1644511149
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1644511149
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1644511149
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_153
timestamp 1644511149
transform 1 0 15180 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_159
timestamp 1644511149
transform 1 0 15732 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_167
timestamp 1644511149
transform 1 0 16468 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_177
timestamp 1644511149
transform 1 0 17388 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_185
timestamp 1644511149
transform 1 0 18124 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_205
timestamp 1644511149
transform 1 0 19964 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_209
timestamp 1644511149
transform 1 0 20332 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_218
timestamp 1644511149
transform 1 0 21160 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_227
timestamp 1644511149
transform 1 0 21988 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_44_272
timestamp 1644511149
transform 1 0 26128 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_294
timestamp 1644511149
transform 1 0 28152 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1644511149
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_317
timestamp 1644511149
transform 1 0 30268 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_324
timestamp 1644511149
transform 1 0 30912 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_328
timestamp 1644511149
transform 1 0 31280 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_337
timestamp 1644511149
transform 1 0 32108 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_341
timestamp 1644511149
transform 1 0 32476 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_348
timestamp 1644511149
transform 1 0 33120 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1644511149
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_373
timestamp 1644511149
transform 1 0 35420 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_384
timestamp 1644511149
transform 1 0 36432 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_392
timestamp 1644511149
transform 1 0 37168 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_397
timestamp 1644511149
transform 1 0 37628 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1644511149
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1644511149
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1644511149
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1644511149
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1644511149
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1644511149
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_73
timestamp 1644511149
transform 1 0 7820 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_83
timestamp 1644511149
transform 1 0 8740 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_95
timestamp 1644511149
transform 1 0 9844 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_107
timestamp 1644511149
transform 1 0 10948 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_137
timestamp 1644511149
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_158
timestamp 1644511149
transform 1 0 15640 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_166
timestamp 1644511149
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_176
timestamp 1644511149
transform 1 0 17296 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_184
timestamp 1644511149
transform 1 0 18032 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_188
timestamp 1644511149
transform 1 0 18400 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_197
timestamp 1644511149
transform 1 0 19228 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_211
timestamp 1644511149
transform 1 0 20516 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_215
timestamp 1644511149
transform 1 0 20884 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1644511149
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_231
timestamp 1644511149
transform 1 0 22356 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_241
timestamp 1644511149
transform 1 0 23276 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_253
timestamp 1644511149
transform 1 0 24380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_265
timestamp 1644511149
transform 1 0 25484 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1644511149
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1644511149
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_289
timestamp 1644511149
transform 1 0 27692 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_313
timestamp 1644511149
transform 1 0 29900 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_321
timestamp 1644511149
transform 1 0 30636 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_333
timestamp 1644511149
transform 1 0 31740 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_383
timestamp 1644511149
transform 1 0 36340 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_401
timestamp 1644511149
transform 1 0 37996 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1644511149
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1644511149
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_71
timestamp 1644511149
transform 1 0 7636 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_76
timestamp 1644511149
transform 1 0 8096 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_85
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_109
timestamp 1644511149
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_121
timestamp 1644511149
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_159
timestamp 1644511149
transform 1 0 15732 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_172
timestamp 1644511149
transform 1 0 16928 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_176
timestamp 1644511149
transform 1 0 17296 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_180
timestamp 1644511149
transform 1 0 17664 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_200
timestamp 1644511149
transform 1 0 19504 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_206
timestamp 1644511149
transform 1 0 20056 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_215
timestamp 1644511149
transform 1 0 20884 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_223
timestamp 1644511149
transform 1 0 21620 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_231
timestamp 1644511149
transform 1 0 22356 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_243
timestamp 1644511149
transform 1 0 23460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1644511149
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_265
timestamp 1644511149
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_277
timestamp 1644511149
transform 1 0 26588 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_289
timestamp 1644511149
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_317
timestamp 1644511149
transform 1 0 30268 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_324
timestamp 1644511149
transform 1 0 30912 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_344
timestamp 1644511149
transform 1 0 32752 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1644511149
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1644511149
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_381
timestamp 1644511149
transform 1 0 36156 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_403
timestamp 1644511149
transform 1 0 38180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1644511149
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_69
timestamp 1644511149
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1644511149
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1644511149
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_132
timestamp 1644511149
transform 1 0 13248 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_148
timestamp 1644511149
transform 1 0 14720 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_164
timestamp 1644511149
transform 1 0 16192 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_175
timestamp 1644511149
transform 1 0 17204 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1644511149
transform 1 0 18032 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_200
timestamp 1644511149
transform 1 0 19504 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_220
timestamp 1644511149
transform 1 0 21344 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_228
timestamp 1644511149
transform 1 0 22080 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_237
timestamp 1644511149
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_249
timestamp 1644511149
transform 1 0 24012 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_253
timestamp 1644511149
transform 1 0 24380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_258
timestamp 1644511149
transform 1 0 24840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_267
timestamp 1644511149
transform 1 0 25668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1644511149
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_285
timestamp 1644511149
transform 1 0 27324 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_298
timestamp 1644511149
transform 1 0 28520 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_306
timestamp 1644511149
transform 1 0 29256 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_318
timestamp 1644511149
transform 1 0 30360 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_326
timestamp 1644511149
transform 1 0 31096 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_343
timestamp 1644511149
transform 1 0 32660 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_348
timestamp 1644511149
transform 1 0 33120 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_359
timestamp 1644511149
transform 1 0 34132 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1644511149
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_396
timestamp 1644511149
transform 1 0 37536 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_403
timestamp 1644511149
transform 1 0 38180 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_14
timestamp 1644511149
transform 1 0 2392 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_26
timestamp 1644511149
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1644511149
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1644511149
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_85
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_109
timestamp 1644511149
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_121
timestamp 1644511149
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1644511149
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1644511149
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_157
timestamp 1644511149
transform 1 0 15548 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_177
timestamp 1644511149
transform 1 0 17388 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_183
timestamp 1644511149
transform 1 0 17940 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_209
timestamp 1644511149
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_221
timestamp 1644511149
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_233
timestamp 1644511149
transform 1 0 22540 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_242
timestamp 1644511149
transform 1 0 23368 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_250
timestamp 1644511149
transform 1 0 24104 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_269
timestamp 1644511149
transform 1 0 25852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_277
timestamp 1644511149
transform 1 0 26588 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_284
timestamp 1644511149
transform 1 0 27232 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_291
timestamp 1644511149
transform 1 0 27876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_295
timestamp 1644511149
transform 1 0 28244 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1644511149
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_321
timestamp 1644511149
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_333
timestamp 1644511149
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_345
timestamp 1644511149
transform 1 0 32844 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_358
timestamp 1644511149
transform 1 0 34040 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_371
timestamp 1644511149
transform 1 0 35236 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_396
timestamp 1644511149
transform 1 0 37536 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_403
timestamp 1644511149
transform 1 0 38180 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1644511149
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1644511149
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_137
timestamp 1644511149
transform 1 0 13708 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_145
timestamp 1644511149
transform 1 0 14444 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1644511149
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1644511149
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_169
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_181
timestamp 1644511149
transform 1 0 17756 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_199
timestamp 1644511149
transform 1 0 19412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_211
timestamp 1644511149
transform 1 0 20516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_231
timestamp 1644511149
transform 1 0 22356 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_249
timestamp 1644511149
transform 1 0 24012 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_257
timestamp 1644511149
transform 1 0 24748 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_262
timestamp 1644511149
transform 1 0 25208 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_274
timestamp 1644511149
transform 1 0 26312 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_297
timestamp 1644511149
transform 1 0 28428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_305
timestamp 1644511149
transform 1 0 29164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_311
timestamp 1644511149
transform 1 0 29716 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_325
timestamp 1644511149
transform 1 0 31004 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_332
timestamp 1644511149
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_358
timestamp 1644511149
transform 1 0 34040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_365
timestamp 1644511149
transform 1 0 34684 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_373
timestamp 1644511149
transform 1 0 35420 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_379
timestamp 1644511149
transform 1 0 35972 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1644511149
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_396
timestamp 1644511149
transform 1 0 37536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_403
timestamp 1644511149
transform 1 0 38180 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_3
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_10
timestamp 1644511149
transform 1 0 2024 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_22
timestamp 1644511149
transform 1 0 3128 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_97
timestamp 1644511149
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_121
timestamp 1644511149
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1644511149
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_146
timestamp 1644511149
transform 1 0 14536 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_166
timestamp 1644511149
transform 1 0 16376 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_178
timestamp 1644511149
transform 1 0 17480 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_190
timestamp 1644511149
transform 1 0 18584 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_209
timestamp 1644511149
transform 1 0 20332 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_219
timestamp 1644511149
transform 1 0 21252 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_229
timestamp 1644511149
transform 1 0 22172 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_237
timestamp 1644511149
transform 1 0 22908 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_243
timestamp 1644511149
transform 1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1644511149
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_261
timestamp 1644511149
transform 1 0 25116 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_266
timestamp 1644511149
transform 1 0 25576 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_273
timestamp 1644511149
transform 1 0 26220 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_279
timestamp 1644511149
transform 1 0 26772 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_283
timestamp 1644511149
transform 1 0 27140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_295
timestamp 1644511149
transform 1 0 28244 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_299
timestamp 1644511149
transform 1 0 28612 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_304
timestamp 1644511149
transform 1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_325
timestamp 1644511149
transform 1 0 31004 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_333
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_341
timestamp 1644511149
transform 1 0 32476 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_348
timestamp 1644511149
transform 1 0 33120 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_360
timestamp 1644511149
transform 1 0 34224 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_370
timestamp 1644511149
transform 1 0 35144 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1644511149
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_81
timestamp 1644511149
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1644511149
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1644511149
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1644511149
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_137
timestamp 1644511149
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_158
timestamp 1644511149
transform 1 0 15640 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_166
timestamp 1644511149
transform 1 0 16376 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_169
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_191
timestamp 1644511149
transform 1 0 18676 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_203
timestamp 1644511149
transform 1 0 19780 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_232
timestamp 1644511149
transform 1 0 22448 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_244
timestamp 1644511149
transform 1 0 23552 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_256
timestamp 1644511149
transform 1 0 24656 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_285
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_289
timestamp 1644511149
transform 1 0 27692 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_297
timestamp 1644511149
transform 1 0 28428 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_304
timestamp 1644511149
transform 1 0 29072 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_311
timestamp 1644511149
transform 1 0 29716 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_315
timestamp 1644511149
transform 1 0 30084 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_345
timestamp 1644511149
transform 1 0 32844 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_354
timestamp 1644511149
transform 1 0 33672 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_374
timestamp 1644511149
transform 1 0 35512 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_382
timestamp 1644511149
transform 1 0 36248 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1644511149
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_397
timestamp 1644511149
transform 1 0 37628 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_109
timestamp 1644511149
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_121
timestamp 1644511149
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1644511149
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1644511149
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_141
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_146
timestamp 1644511149
transform 1 0 14536 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_166
timestamp 1644511149
transform 1 0 16376 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_186
timestamp 1644511149
transform 1 0 18216 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1644511149
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_197
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_203
timestamp 1644511149
transform 1 0 19780 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_209
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_219
timestamp 1644511149
transform 1 0 21252 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_226
timestamp 1644511149
transform 1 0 21896 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_242
timestamp 1644511149
transform 1 0 23368 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1644511149
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_259
timestamp 1644511149
transform 1 0 24932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_270
timestamp 1644511149
transform 1 0 25944 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_289
timestamp 1644511149
transform 1 0 27692 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_299
timestamp 1644511149
transform 1 0 28612 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_313
timestamp 1644511149
transform 1 0 29900 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_320
timestamp 1644511149
transform 1 0 30544 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_332
timestamp 1644511149
transform 1 0 31648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_346
timestamp 1644511149
transform 1 0 32936 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_358
timestamp 1644511149
transform 1 0 34040 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_381
timestamp 1644511149
transform 1 0 36156 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1644511149
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1644511149
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1644511149
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1644511149
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1644511149
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_137
timestamp 1644511149
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_149
timestamp 1644511149
transform 1 0 14812 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_53_160
timestamp 1644511149
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_174
timestamp 1644511149
transform 1 0 17112 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_187
timestamp 1644511149
transform 1 0 18308 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_204
timestamp 1644511149
transform 1 0 19872 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_210
timestamp 1644511149
transform 1 0 20424 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_219
timestamp 1644511149
transform 1 0 21252 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1644511149
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_233
timestamp 1644511149
transform 1 0 22540 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_251
timestamp 1644511149
transform 1 0 24196 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_257
timestamp 1644511149
transform 1 0 24748 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_265
timestamp 1644511149
transform 1 0 25484 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_276
timestamp 1644511149
transform 1 0 26496 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_281
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_285
timestamp 1644511149
transform 1 0 27324 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_302
timestamp 1644511149
transform 1 0 28888 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_316
timestamp 1644511149
transform 1 0 30176 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_323
timestamp 1644511149
transform 1 0 30820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_353
timestamp 1644511149
transform 1 0 33580 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_365
timestamp 1644511149
transform 1 0 34684 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_371
timestamp 1644511149
transform 1 0 35236 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_388
timestamp 1644511149
transform 1 0 36800 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_398
timestamp 1644511149
transform 1 0 37720 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_406
timestamp 1644511149
transform 1 0 38456 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1644511149
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1644511149
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1644511149
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1644511149
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_97
timestamp 1644511149
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_109
timestamp 1644511149
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_121
timestamp 1644511149
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1644511149
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1644511149
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_147
timestamp 1644511149
transform 1 0 14628 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_151
timestamp 1644511149
transform 1 0 14996 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_160
timestamp 1644511149
transform 1 0 15824 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_166
timestamp 1644511149
transform 1 0 16376 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_173
timestamp 1644511149
transform 1 0 17020 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_181
timestamp 1644511149
transform 1 0 17756 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1644511149
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_201
timestamp 1644511149
transform 1 0 19596 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_218
timestamp 1644511149
transform 1 0 21160 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_230
timestamp 1644511149
transform 1 0 22264 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_236
timestamp 1644511149
transform 1 0 22816 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_241
timestamp 1644511149
transform 1 0 23276 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_249
timestamp 1644511149
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_259
timestamp 1644511149
transform 1 0 24932 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_286
timestamp 1644511149
transform 1 0 27416 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_298
timestamp 1644511149
transform 1 0 28520 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1644511149
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_318
timestamp 1644511149
transform 1 0 30360 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_328
timestamp 1644511149
transform 1 0 31280 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_334
timestamp 1644511149
transform 1 0 31832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_338
timestamp 1644511149
transform 1 0 32200 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_351
timestamp 1644511149
transform 1 0 33396 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_358
timestamp 1644511149
transform 1 0 34040 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_373
timestamp 1644511149
transform 1 0 35420 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_378
timestamp 1644511149
transform 1 0 35880 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_403
timestamp 1644511149
transform 1 0 38180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_137
timestamp 1644511149
transform 1 0 13708 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_159
timestamp 1644511149
transform 1 0 15732 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_176
timestamp 1644511149
transform 1 0 17296 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_184
timestamp 1644511149
transform 1 0 18032 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_202
timestamp 1644511149
transform 1 0 19688 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_213
timestamp 1644511149
transform 1 0 20700 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_221
timestamp 1644511149
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_244
timestamp 1644511149
transform 1 0 23552 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_254
timestamp 1644511149
transform 1 0 24472 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_262
timestamp 1644511149
transform 1 0 25208 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_269
timestamp 1644511149
transform 1 0 25852 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_277
timestamp 1644511149
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_289
timestamp 1644511149
transform 1 0 27692 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_299
timestamp 1644511149
transform 1 0 28612 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_311
timestamp 1644511149
transform 1 0 29716 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_55_322
timestamp 1644511149
transform 1 0 30728 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_332
timestamp 1644511149
transform 1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_343
timestamp 1644511149
transform 1 0 32660 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_363
timestamp 1644511149
transform 1 0 34500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_374
timestamp 1644511149
transform 1 0 35512 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_383
timestamp 1644511149
transform 1 0 36340 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_398
timestamp 1644511149
transform 1 0 37720 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_406
timestamp 1644511149
transform 1 0 38456 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1644511149
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1644511149
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1644511149
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_160
timestamp 1644511149
transform 1 0 15824 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_172
timestamp 1644511149
transform 1 0 16928 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_179
timestamp 1644511149
transform 1 0 17572 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_188
timestamp 1644511149
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_221
timestamp 1644511149
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_233
timestamp 1644511149
transform 1 0 22540 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_241
timestamp 1644511149
transform 1 0 23276 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_247
timestamp 1644511149
transform 1 0 23828 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1644511149
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_277
timestamp 1644511149
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_289
timestamp 1644511149
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1644511149
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1644511149
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_315
timestamp 1644511149
transform 1 0 30084 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_326
timestamp 1644511149
transform 1 0 31096 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_334
timestamp 1644511149
transform 1 0 31832 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_341
timestamp 1644511149
transform 1 0 32476 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_348
timestamp 1644511149
transform 1 0 33120 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1644511149
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_375
timestamp 1644511149
transform 1 0 35604 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_397
timestamp 1644511149
transform 1 0 37628 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1644511149
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1644511149
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1644511149
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1644511149
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1644511149
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_156
timestamp 1644511149
transform 1 0 15456 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_187
timestamp 1644511149
transform 1 0 18308 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_199
timestamp 1644511149
transform 1 0 19412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_211
timestamp 1644511149
transform 1 0 20516 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_215
timestamp 1644511149
transform 1 0 20884 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1644511149
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_229
timestamp 1644511149
transform 1 0 22172 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_241
timestamp 1644511149
transform 1 0 23276 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_253
timestamp 1644511149
transform 1 0 24380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_259
timestamp 1644511149
transform 1 0 24932 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_276
timestamp 1644511149
transform 1 0 26496 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_288
timestamp 1644511149
transform 1 0 27600 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_300
timestamp 1644511149
transform 1 0 28704 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_57_312
timestamp 1644511149
transform 1 0 29808 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_322
timestamp 1644511149
transform 1 0 30728 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_334
timestamp 1644511149
transform 1 0 31832 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_357
timestamp 1644511149
transform 1 0 33948 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_366
timestamp 1644511149
transform 1 0 34776 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_378
timestamp 1644511149
transform 1 0 35880 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_387
timestamp 1644511149
transform 1 0 36708 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1644511149
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_399
timestamp 1644511149
transform 1 0 37812 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_165
timestamp 1644511149
transform 1 0 16284 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_174
timestamp 1644511149
transform 1 0 17112 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1644511149
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1644511149
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_200
timestamp 1644511149
transform 1 0 19504 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_204
timestamp 1644511149
transform 1 0 19872 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_221
timestamp 1644511149
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_233
timestamp 1644511149
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1644511149
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1644511149
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_259
timestamp 1644511149
transform 1 0 24932 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_271
timestamp 1644511149
transform 1 0 26036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_277
timestamp 1644511149
transform 1 0 26588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_286
timestamp 1644511149
transform 1 0 27416 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_290
timestamp 1644511149
transform 1 0 27784 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_297
timestamp 1644511149
transform 1 0 28428 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_305
timestamp 1644511149
transform 1 0 29164 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_316
timestamp 1644511149
transform 1 0 30176 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_324
timestamp 1644511149
transform 1 0 30912 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_330
timestamp 1644511149
transform 1 0 31464 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_341
timestamp 1644511149
transform 1 0 32476 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_349
timestamp 1644511149
transform 1 0 33212 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_360
timestamp 1644511149
transform 1 0 34224 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_370
timestamp 1644511149
transform 1 0 35144 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_383
timestamp 1644511149
transform 1 0 36340 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_403
timestamp 1644511149
transform 1 0 38180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_113
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_125
timestamp 1644511149
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_137
timestamp 1644511149
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_149
timestamp 1644511149
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_188
timestamp 1644511149
transform 1 0 18400 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_208
timestamp 1644511149
transform 1 0 20240 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_219
timestamp 1644511149
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1644511149
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_239
timestamp 1644511149
transform 1 0 23092 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_246
timestamp 1644511149
transform 1 0 23736 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_263
timestamp 1644511149
transform 1 0 25300 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_271
timestamp 1644511149
transform 1 0 26036 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_287
timestamp 1644511149
transform 1 0 27508 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_299
timestamp 1644511149
transform 1 0 28612 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_310
timestamp 1644511149
transform 1 0 29624 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_330
timestamp 1644511149
transform 1 0 31464 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_353
timestamp 1644511149
transform 1 0 33580 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_367
timestamp 1644511149
transform 1 0 34868 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_377
timestamp 1644511149
transform 1 0 35788 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_386
timestamp 1644511149
transform 1 0 36616 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_397
timestamp 1644511149
transform 1 0 37628 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_121
timestamp 1644511149
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_173
timestamp 1644511149
transform 1 0 17020 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_182
timestamp 1644511149
transform 1 0 17848 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_191
timestamp 1644511149
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1644511149
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_215
timestamp 1644511149
transform 1 0 20884 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_227
timestamp 1644511149
transform 1 0 21988 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_238
timestamp 1644511149
transform 1 0 23000 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1644511149
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_262
timestamp 1644511149
transform 1 0 25208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_273
timestamp 1644511149
transform 1 0 26220 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_277
timestamp 1644511149
transform 1 0 26588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_285
timestamp 1644511149
transform 1 0 27324 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_296
timestamp 1644511149
transform 1 0 28336 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_317
timestamp 1644511149
transform 1 0 30268 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_329
timestamp 1644511149
transform 1 0 31372 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_339
timestamp 1644511149
transform 1 0 32292 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_343
timestamp 1644511149
transform 1 0 32660 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_360
timestamp 1644511149
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_381
timestamp 1644511149
transform 1 0 36156 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_390
timestamp 1644511149
transform 1 0 36984 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_399
timestamp 1644511149
transform 1 0 37812 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_12
timestamp 1644511149
transform 1 0 2208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_16
timestamp 1644511149
transform 1 0 2576 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_20
timestamp 1644511149
transform 1 0 2944 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_32
timestamp 1644511149
transform 1 0 4048 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_44
timestamp 1644511149
transform 1 0 5152 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_81
timestamp 1644511149
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_93
timestamp 1644511149
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1644511149
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1644511149
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_178
timestamp 1644511149
transform 1 0 17480 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_190
timestamp 1644511149
transform 1 0 18584 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_202
timestamp 1644511149
transform 1 0 19688 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1644511149
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_244
timestamp 1644511149
transform 1 0 23552 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_252
timestamp 1644511149
transform 1 0 24288 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_261
timestamp 1644511149
transform 1 0 25116 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_268
timestamp 1644511149
transform 1 0 25760 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_289
timestamp 1644511149
transform 1 0 27692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_301
timestamp 1644511149
transform 1 0 28796 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_313
timestamp 1644511149
transform 1 0 29900 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_325
timestamp 1644511149
transform 1 0 31004 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp 1644511149
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_352
timestamp 1644511149
transform 1 0 33488 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_368
timestamp 1644511149
transform 1 0 34960 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_376
timestamp 1644511149
transform 1 0 35696 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_382
timestamp 1644511149
transform 1 0 36248 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1644511149
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1644511149
transform 1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_24
timestamp 1644511149
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_65
timestamp 1644511149
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1644511149
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1644511149
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_146
timestamp 1644511149
transform 1 0 14536 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_158
timestamp 1644511149
transform 1 0 15640 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_170
timestamp 1644511149
transform 1 0 16744 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_182
timestamp 1644511149
transform 1 0 17848 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_194
timestamp 1644511149
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_197
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_205
timestamp 1644511149
transform 1 0 19964 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_211
timestamp 1644511149
transform 1 0 20516 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_219
timestamp 1644511149
transform 1 0 21252 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_225
timestamp 1644511149
transform 1 0 21804 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_237
timestamp 1644511149
transform 1 0 22908 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1644511149
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_257
timestamp 1644511149
transform 1 0 24748 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_265
timestamp 1644511149
transform 1 0 25484 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_272
timestamp 1644511149
transform 1 0 26128 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_280
timestamp 1644511149
transform 1 0 26864 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_286
timestamp 1644511149
transform 1 0 27416 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_298
timestamp 1644511149
transform 1 0 28520 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_306
timestamp 1644511149
transform 1 0 29256 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_332
timestamp 1644511149
transform 1 0 31648 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_344
timestamp 1644511149
transform 1 0 32752 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_356
timestamp 1644511149
transform 1 0 33856 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_381
timestamp 1644511149
transform 1 0 36156 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_398
timestamp 1644511149
transform 1 0 37720 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1644511149
transform 1 0 38456 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1644511149
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1644511149
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1644511149
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1644511149
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1644511149
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_69
timestamp 1644511149
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_81
timestamp 1644511149
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_93
timestamp 1644511149
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1644511149
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1644511149
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_189
timestamp 1644511149
transform 1 0 18492 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_206
timestamp 1644511149
transform 1 0 20056 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_218
timestamp 1644511149
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_233
timestamp 1644511149
transform 1 0 22540 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_240
timestamp 1644511149
transform 1 0 23184 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_247
timestamp 1644511149
transform 1 0 23828 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_259
timestamp 1644511149
transform 1 0 24932 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_63_266
timestamp 1644511149
transform 1 0 25576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_274
timestamp 1644511149
transform 1 0 26312 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_281
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_288
timestamp 1644511149
transform 1 0 27600 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_300
timestamp 1644511149
transform 1 0 28704 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_308
timestamp 1644511149
transform 1 0 29440 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_315
timestamp 1644511149
transform 1 0 30084 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_323
timestamp 1644511149
transform 1 0 30820 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1644511149
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1644511149
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_353
timestamp 1644511149
transform 1 0 33580 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_388
timestamp 1644511149
transform 1 0 36800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_397
timestamp 1644511149
transform 1 0 37628 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1644511149
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1644511149
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_160
timestamp 1644511149
transform 1 0 15824 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_168
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_173
timestamp 1644511149
transform 1 0 17020 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_177
timestamp 1644511149
transform 1 0 17388 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_185
timestamp 1644511149
transform 1 0 18124 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1644511149
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_202
timestamp 1644511149
transform 1 0 19688 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_210
timestamp 1644511149
transform 1 0 20424 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_227
timestamp 1644511149
transform 1 0 21988 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_239
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_256
timestamp 1644511149
transform 1 0 24656 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_274
timestamp 1644511149
transform 1 0 26312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_285
timestamp 1644511149
transform 1 0 27324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_292
timestamp 1644511149
transform 1 0 27968 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_296
timestamp 1644511149
transform 1 0 28336 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1644511149
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_325
timestamp 1644511149
transform 1 0 31004 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_331
timestamp 1644511149
transform 1 0 31556 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_341
timestamp 1644511149
transform 1 0 32476 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_350
timestamp 1644511149
transform 1 0 33304 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_362
timestamp 1644511149
transform 1 0 34408 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_370
timestamp 1644511149
transform 1 0 35144 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_374
timestamp 1644511149
transform 1 0 35512 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_378
timestamp 1644511149
transform 1 0 35880 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1644511149
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1644511149
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1644511149
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1644511149
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1644511149
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_144
timestamp 1644511149
transform 1 0 14352 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_156
timestamp 1644511149
transform 1 0 15456 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_160
timestamp 1644511149
transform 1 0 15824 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_164
timestamp 1644511149
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_185
timestamp 1644511149
transform 1 0 18124 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_194
timestamp 1644511149
transform 1 0 18952 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_201
timestamp 1644511149
transform 1 0 19596 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_205
timestamp 1644511149
transform 1 0 19964 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_213
timestamp 1644511149
transform 1 0 20700 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_237
timestamp 1644511149
transform 1 0 22908 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_242
timestamp 1644511149
transform 1 0 23368 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_252
timestamp 1644511149
transform 1 0 24288 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_260
timestamp 1644511149
transform 1 0 25024 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_268
timestamp 1644511149
transform 1 0 25760 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_276
timestamp 1644511149
transform 1 0 26496 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_289
timestamp 1644511149
transform 1 0 27692 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_65_297
timestamp 1644511149
transform 1 0 28428 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_307
timestamp 1644511149
transform 1 0 29348 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_315
timestamp 1644511149
transform 1 0 30084 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_327
timestamp 1644511149
transform 1 0 31188 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1644511149
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_346
timestamp 1644511149
transform 1 0 32936 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_358
timestamp 1644511149
transform 1 0 34040 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_364
timestamp 1644511149
transform 1 0 34592 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_65_388
timestamp 1644511149
transform 1 0 36800 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_397
timestamp 1644511149
transform 1 0 37628 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_7
timestamp 1644511149
transform 1 0 1748 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_11
timestamp 1644511149
transform 1 0 2116 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_66_20
timestamp 1644511149
transform 1 0 2944 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_172
timestamp 1644511149
transform 1 0 16928 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_178
timestamp 1644511149
transform 1 0 17480 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_185
timestamp 1644511149
transform 1 0 18124 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_193
timestamp 1644511149
transform 1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_203
timestamp 1644511149
transform 1 0 19780 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_210
timestamp 1644511149
transform 1 0 20424 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_219
timestamp 1644511149
transform 1 0 21252 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_227
timestamp 1644511149
transform 1 0 21988 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_66_246
timestamp 1644511149
transform 1 0 23736 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_260
timestamp 1644511149
transform 1 0 25024 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_272
timestamp 1644511149
transform 1 0 26128 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_284
timestamp 1644511149
transform 1 0 27232 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_302
timestamp 1644511149
transform 1 0 28888 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_309
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_321
timestamp 1644511149
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_333
timestamp 1644511149
transform 1 0 31740 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_345
timestamp 1644511149
transform 1 0 32844 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_354
timestamp 1644511149
transform 1 0 33672 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_362
timestamp 1644511149
transform 1 0 34408 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_378
timestamp 1644511149
transform 1 0 35880 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_403
timestamp 1644511149
transform 1 0 38180 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_7
timestamp 1644511149
transform 1 0 1748 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_29
timestamp 1644511149
transform 1 0 3772 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_41
timestamp 1644511149
transform 1 0 4876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_53
timestamp 1644511149
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_146
timestamp 1644511149
transform 1 0 14536 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_158
timestamp 1644511149
transform 1 0 15640 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_166
timestamp 1644511149
transform 1 0 16376 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_174
timestamp 1644511149
transform 1 0 17112 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_186
timestamp 1644511149
transform 1 0 18216 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_192
timestamp 1644511149
transform 1 0 18768 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_204
timestamp 1644511149
transform 1 0 19872 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_210
timestamp 1644511149
transform 1 0 20424 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_230
timestamp 1644511149
transform 1 0 22264 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_242
timestamp 1644511149
transform 1 0 23368 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_254
timestamp 1644511149
transform 1 0 24472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_264
timestamp 1644511149
transform 1 0 25392 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_274
timestamp 1644511149
transform 1 0 26312 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1644511149
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_305
timestamp 1644511149
transform 1 0 29164 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_313
timestamp 1644511149
transform 1 0 29900 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_332
timestamp 1644511149
transform 1 0 31648 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_342
timestamp 1644511149
transform 1 0 32568 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_354
timestamp 1644511149
transform 1 0 33672 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_366
timestamp 1644511149
transform 1 0 34776 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_67_388
timestamp 1644511149
transform 1 0 36800 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_398
timestamp 1644511149
transform 1 0 37720 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_406
timestamp 1644511149
transform 1 0 38456 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_12
timestamp 1644511149
transform 1 0 2208 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_24
timestamp 1644511149
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_169
timestamp 1644511149
transform 1 0 16652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_175
timestamp 1644511149
transform 1 0 17204 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_186
timestamp 1644511149
transform 1 0 18216 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_194
timestamp 1644511149
transform 1 0 18952 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_197
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_68_219
timestamp 1644511149
transform 1 0 21252 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_227
timestamp 1644511149
transform 1 0 21988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_239
timestamp 1644511149
transform 1 0 23092 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1644511149
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_253
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_264
timestamp 1644511149
transform 1 0 25392 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_276
timestamp 1644511149
transform 1 0 26496 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_288
timestamp 1644511149
transform 1 0 27600 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_68_299
timestamp 1644511149
transform 1 0 28612 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1644511149
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_321
timestamp 1644511149
transform 1 0 30636 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_327
timestamp 1644511149
transform 1 0 31188 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_335
timestamp 1644511149
transform 1 0 31924 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_341
timestamp 1644511149
transform 1 0 32476 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_348
timestamp 1644511149
transform 1 0 33120 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_356
timestamp 1644511149
transform 1 0 33856 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_360
timestamp 1644511149
transform 1 0 34224 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_68_372
timestamp 1644511149
transform 1 0 35328 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_380
timestamp 1644511149
transform 1 0 36064 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_403
timestamp 1644511149
transform 1 0 38180 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_26
timestamp 1644511149
transform 1 0 3496 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_38
timestamp 1644511149
transform 1 0 4600 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_50
timestamp 1644511149
transform 1 0 5704 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_185
timestamp 1644511149
transform 1 0 18124 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_205
timestamp 1644511149
transform 1 0 19964 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_214
timestamp 1644511149
transform 1 0 20792 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_222
timestamp 1644511149
transform 1 0 21528 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_235
timestamp 1644511149
transform 1 0 22724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_247
timestamp 1644511149
transform 1 0 23828 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_69_255
timestamp 1644511149
transform 1 0 24564 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_262
timestamp 1644511149
transform 1 0 25208 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_269
timestamp 1644511149
transform 1 0 25852 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_277
timestamp 1644511149
transform 1 0 26588 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_286
timestamp 1644511149
transform 1 0 27416 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_298
timestamp 1644511149
transform 1 0 28520 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_69_317
timestamp 1644511149
transform 1 0 30268 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_325
timestamp 1644511149
transform 1 0 31004 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_332
timestamp 1644511149
transform 1 0 31648 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_353
timestamp 1644511149
transform 1 0 33580 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_382
timestamp 1644511149
transform 1 0 36248 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_390
timestamp 1644511149
transform 1 0 36984 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_396
timestamp 1644511149
transform 1 0 37536 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_403
timestamp 1644511149
transform 1 0 38180 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_8
timestamp 1644511149
transform 1 0 1840 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_20
timestamp 1644511149
transform 1 0 2944 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_113
timestamp 1644511149
transform 1 0 11500 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_125
timestamp 1644511149
transform 1 0 12604 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_137
timestamp 1644511149
transform 1 0 13708 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_170
timestamp 1644511149
transform 1 0 16744 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_182
timestamp 1644511149
transform 1 0 17848 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_194
timestamp 1644511149
transform 1 0 18952 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_207
timestamp 1644511149
transform 1 0 20148 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_70_219
timestamp 1644511149
transform 1 0 21252 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_239
timestamp 1644511149
transform 1 0 23092 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_248
timestamp 1644511149
transform 1 0 23920 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_262
timestamp 1644511149
transform 1 0 25208 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_272
timestamp 1644511149
transform 1 0 26128 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_276
timestamp 1644511149
transform 1 0 26496 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_293
timestamp 1644511149
transform 1 0 28060 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_305
timestamp 1644511149
transform 1 0 29164 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_341
timestamp 1644511149
transform 1 0 32476 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_346
timestamp 1644511149
transform 1 0 32936 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_354
timestamp 1644511149
transform 1 0 33672 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_360
timestamp 1644511149
transform 1 0 34224 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_371
timestamp 1644511149
transform 1 0 35236 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_378
timestamp 1644511149
transform 1 0 35880 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_403
timestamp 1644511149
transform 1 0 38180 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1644511149
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1644511149
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_51
timestamp 1644511149
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1644511149
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_77
timestamp 1644511149
transform 1 0 8188 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_84
timestamp 1644511149
transform 1 0 8832 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_108
timestamp 1644511149
transform 1 0 11040 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_203
timestamp 1644511149
transform 1 0 19780 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_215
timestamp 1644511149
transform 1 0 20884 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_225
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_233
timestamp 1644511149
transform 1 0 22540 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_250
timestamp 1644511149
transform 1 0 24104 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_256
timestamp 1644511149
transform 1 0 24656 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_262
timestamp 1644511149
transform 1 0 25208 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_274
timestamp 1644511149
transform 1 0 26312 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_284
timestamp 1644511149
transform 1 0 27232 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_296
timestamp 1644511149
transform 1 0 28336 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_315
timestamp 1644511149
transform 1 0 30084 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_323
timestamp 1644511149
transform 1 0 30820 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_327
timestamp 1644511149
transform 1 0 31188 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_356
timestamp 1644511149
transform 1 0 33856 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_365
timestamp 1644511149
transform 1 0 34684 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_374
timestamp 1644511149
transform 1 0 35512 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_381
timestamp 1644511149
transform 1 0 36156 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_388
timestamp 1644511149
transform 1 0 36800 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_397
timestamp 1644511149
transform 1 0 37628 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_7
timestamp 1644511149
transform 1 0 1748 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_15
timestamp 1644511149
transform 1 0 2484 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_72_21
timestamp 1644511149
transform 1 0 3036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1644511149
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_105
timestamp 1644511149
transform 1 0 10764 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_117
timestamp 1644511149
transform 1 0 11868 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_129
timestamp 1644511149
transform 1 0 12972 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_137
timestamp 1644511149
transform 1 0 13708 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_161
timestamp 1644511149
transform 1 0 15916 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_72_180
timestamp 1644511149
transform 1 0 17664 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_191
timestamp 1644511149
transform 1 0 18676 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_197
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_203
timestamp 1644511149
transform 1 0 19780 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_209
timestamp 1644511149
transform 1 0 20332 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_216
timestamp 1644511149
transform 1 0 20976 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_228
timestamp 1644511149
transform 1 0 22080 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_234
timestamp 1644511149
transform 1 0 22632 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_238
timestamp 1644511149
transform 1 0 23000 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_250
timestamp 1644511149
transform 1 0 24104 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_273
timestamp 1644511149
transform 1 0 26220 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_290
timestamp 1644511149
transform 1 0 27784 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_298
timestamp 1644511149
transform 1 0 28520 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_304
timestamp 1644511149
transform 1 0 29072 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_314
timestamp 1644511149
transform 1 0 29992 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_322
timestamp 1644511149
transform 1 0 30728 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_326
timestamp 1644511149
transform 1 0 31096 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_351
timestamp 1644511149
transform 1 0 33396 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_360
timestamp 1644511149
transform 1 0 34224 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_381
timestamp 1644511149
transform 1 0 36156 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_403
timestamp 1644511149
transform 1 0 38180 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_6
timestamp 1644511149
transform 1 0 1656 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_31
timestamp 1644511149
transform 1 0 3956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_43
timestamp 1644511149
transform 1 0 5060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_89
timestamp 1644511149
transform 1 0 9292 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_104
timestamp 1644511149
transform 1 0 10672 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_200
timestamp 1644511149
transform 1 0 19504 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_220
timestamp 1644511149
transform 1 0 21344 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_236
timestamp 1644511149
transform 1 0 22816 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_244
timestamp 1644511149
transform 1 0 23552 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_249
timestamp 1644511149
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_261
timestamp 1644511149
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1644511149
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_289
timestamp 1644511149
transform 1 0 27692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_301
timestamp 1644511149
transform 1 0 28796 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_73_313
timestamp 1644511149
transform 1 0 29900 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_323
timestamp 1644511149
transform 1 0 30820 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_369
timestamp 1644511149
transform 1 0 35052 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_381
timestamp 1644511149
transform 1 0 36156 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_388
timestamp 1644511149
transform 1 0 36800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_398
timestamp 1644511149
transform 1 0 37720 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_406
timestamp 1644511149
transform 1 0 38456 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_24
timestamp 1644511149
transform 1 0 3312 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_74_161
timestamp 1644511149
transform 1 0 15916 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_74_167
timestamp 1644511149
transform 1 0 16468 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_176
timestamp 1644511149
transform 1 0 17296 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_188
timestamp 1644511149
transform 1 0 18400 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_192
timestamp 1644511149
transform 1 0 18768 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_74_212
timestamp 1644511149
transform 1 0 20608 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_228
timestamp 1644511149
transform 1 0 22080 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_74_237
timestamp 1644511149
transform 1 0 22908 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_248
timestamp 1644511149
transform 1 0 23920 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_257
timestamp 1644511149
transform 1 0 24748 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_274
timestamp 1644511149
transform 1 0 26312 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_278
timestamp 1644511149
transform 1 0 26680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_285
timestamp 1644511149
transform 1 0 27324 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_294
timestamp 1644511149
transform 1 0 28152 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_306
timestamp 1644511149
transform 1 0 29256 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_316
timestamp 1644511149
transform 1 0 30176 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_322
timestamp 1644511149
transform 1 0 30728 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_339
timestamp 1644511149
transform 1 0 32292 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_351
timestamp 1644511149
transform 1 0 33396 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_381
timestamp 1644511149
transform 1 0 36156 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_403
timestamp 1644511149
transform 1 0 38180 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_8
timestamp 1644511149
transform 1 0 1840 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_186
timestamp 1644511149
transform 1 0 18216 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_194
timestamp 1644511149
transform 1 0 18952 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_200
timestamp 1644511149
transform 1 0 19504 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_210
timestamp 1644511149
transform 1 0 20424 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_222
timestamp 1644511149
transform 1 0 21528 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_233
timestamp 1644511149
transform 1 0 22540 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_244
timestamp 1644511149
transform 1 0 23552 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_264
timestamp 1644511149
transform 1 0 25392 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_288
timestamp 1644511149
transform 1 0 27600 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_300
timestamp 1644511149
transform 1 0 28704 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_308
timestamp 1644511149
transform 1 0 29440 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_314
timestamp 1644511149
transform 1 0 29992 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_377
timestamp 1644511149
transform 1 0 35788 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_381
timestamp 1644511149
transform 1 0 36156 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_388
timestamp 1644511149
transform 1 0 36800 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_397
timestamp 1644511149
transform 1 0 37628 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1644511149
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_27
timestamp 1644511149
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_171
timestamp 1644511149
transform 1 0 16836 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_178
timestamp 1644511149
transform 1 0 17480 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_190
timestamp 1644511149
transform 1 0 18584 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_200
timestamp 1644511149
transform 1 0 19504 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_212
timestamp 1644511149
transform 1 0 20608 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_220
timestamp 1644511149
transform 1 0 21344 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_228
timestamp 1644511149
transform 1 0 22080 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_240
timestamp 1644511149
transform 1 0 23184 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_264
timestamp 1644511149
transform 1 0 25392 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_271
timestamp 1644511149
transform 1 0 26036 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_76_284
timestamp 1644511149
transform 1 0 27232 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_304
timestamp 1644511149
transform 1 0 29072 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_325
timestamp 1644511149
transform 1 0 31004 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_337
timestamp 1644511149
transform 1 0 32108 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_349
timestamp 1644511149
transform 1 0 33212 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_361
timestamp 1644511149
transform 1 0 34316 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_381
timestamp 1644511149
transform 1 0 36156 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_403
timestamp 1644511149
transform 1 0 38180 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1644511149
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_201
timestamp 1644511149
transform 1 0 19596 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_77_208
timestamp 1644511149
transform 1 0 20240 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_77_219
timestamp 1644511149
transform 1 0 21252 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_245
timestamp 1644511149
transform 1 0 23644 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_257
timestamp 1644511149
transform 1 0 24748 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_274
timestamp 1644511149
transform 1 0 26312 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_77_284
timestamp 1644511149
transform 1 0 27232 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_77_314
timestamp 1644511149
transform 1 0 29992 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_326
timestamp 1644511149
transform 1 0 31096 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_334
timestamp 1644511149
transform 1 0 31832 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_388
timestamp 1644511149
transform 1 0 36800 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_397
timestamp 1644511149
transform 1 0 37628 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_8
timestamp 1644511149
transform 1 0 1840 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1644511149
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1644511149
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_78_62
timestamp 1644511149
transform 1 0 6808 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_69
timestamp 1644511149
transform 1 0 7452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_78_81
timestamp 1644511149
transform 1 0 8556 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_78_205
timestamp 1644511149
transform 1 0 19964 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_213
timestamp 1644511149
transform 1 0 20700 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_230
timestamp 1644511149
transform 1 0 22264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_241
timestamp 1644511149
transform 1 0 23276 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_248
timestamp 1644511149
transform 1 0 23920 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_258
timestamp 1644511149
transform 1 0 24840 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_262
timestamp 1644511149
transform 1 0 25208 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_279
timestamp 1644511149
transform 1 0 26772 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_288
timestamp 1644511149
transform 1 0 27600 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_300
timestamp 1644511149
transform 1 0 28704 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_381
timestamp 1644511149
transform 1 0 36156 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_403
timestamp 1644511149
transform 1 0 38180 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_13
timestamp 1644511149
transform 1 0 2300 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_20
timestamp 1644511149
transform 1 0 2944 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1644511149
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_39
timestamp 1644511149
transform 1 0 4692 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_47
timestamp 1644511149
transform 1 0 5428 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_52
timestamp 1644511149
transform 1 0 5888 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_80
timestamp 1644511149
transform 1 0 8464 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_87
timestamp 1644511149
transform 1 0 9108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_99
timestamp 1644511149
transform 1 0 10212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_155
timestamp 1644511149
transform 1 0 15364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_177
timestamp 1644511149
transform 1 0 17388 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_199
timestamp 1644511149
transform 1 0 19412 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_219
timestamp 1644511149
transform 1 0 21252 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_235
timestamp 1644511149
transform 1 0 22724 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_259
timestamp 1644511149
transform 1 0 24932 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_266
timestamp 1644511149
transform 1 0 25576 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_272
timestamp 1644511149
transform 1 0 26128 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_276
timestamp 1644511149
transform 1 0 26496 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_297
timestamp 1644511149
transform 1 0 28428 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_308
timestamp 1644511149
transform 1 0 29440 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_320
timestamp 1644511149
transform 1 0 30544 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_324
timestamp 1644511149
transform 1 0 30912 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_328
timestamp 1644511149
transform 1 0 31280 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_340
timestamp 1644511149
transform 1 0 32384 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_352
timestamp 1644511149
transform 1 0 33488 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_364
timestamp 1644511149
transform 1 0 34592 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_388
timestamp 1644511149
transform 1 0 36800 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_396
timestamp 1644511149
transform 1 0 37536 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_403
timestamp 1644511149
transform 1 0 38180 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_24
timestamp 1644511149
transform 1 0 3312 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_32
timestamp 1644511149
transform 1 0 4048 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_36
timestamp 1644511149
transform 1 0 4416 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_40
timestamp 1644511149
transform 1 0 4784 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_47
timestamp 1644511149
transform 1 0 5428 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_72
timestamp 1644511149
transform 1 0 7728 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_79
timestamp 1644511149
transform 1 0 8372 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1644511149
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_106
timestamp 1644511149
transform 1 0 10856 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_118
timestamp 1644511149
transform 1 0 11960 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_130
timestamp 1644511149
transform 1 0 13064 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_138
timestamp 1644511149
transform 1 0 13800 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_149
timestamp 1644511149
transform 1 0 14812 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_171
timestamp 1644511149
transform 1 0 16836 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_178
timestamp 1644511149
transform 1 0 17480 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_184
timestamp 1644511149
transform 1 0 18032 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_188
timestamp 1644511149
transform 1 0 18400 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_80_200
timestamp 1644511149
transform 1 0 19504 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_206
timestamp 1644511149
transform 1 0 20056 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_228
timestamp 1644511149
transform 1 0 22080 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_235
timestamp 1644511149
transform 1 0 22724 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_247
timestamp 1644511149
transform 1 0 23828 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_256
timestamp 1644511149
transform 1 0 24656 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_268
timestamp 1644511149
transform 1 0 25760 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_272
timestamp 1644511149
transform 1 0 26128 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_294
timestamp 1644511149
transform 1 0 28152 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1644511149
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_312
timestamp 1644511149
transform 1 0 29808 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_352
timestamp 1644511149
transform 1 0 33488 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_359
timestamp 1644511149
transform 1 0 34132 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_381
timestamp 1644511149
transform 1 0 36156 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_403
timestamp 1644511149
transform 1 0 38180 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_6
timestamp 1644511149
transform 1 0 1656 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_31
timestamp 1644511149
transform 1 0 3956 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_45
timestamp 1644511149
transform 1 0 5244 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_52
timestamp 1644511149
transform 1 0 5888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_60
timestamp 1644511149
transform 1 0 6624 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_66
timestamp 1644511149
transform 1 0 7176 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_70
timestamp 1644511149
transform 1 0 7544 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_95
timestamp 1644511149
transform 1 0 9844 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_107
timestamp 1644511149
transform 1 0 10948 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_81_154
timestamp 1644511149
transform 1 0 15272 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_160
timestamp 1644511149
transform 1 0 15824 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_164
timestamp 1644511149
transform 1 0 16192 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_173
timestamp 1644511149
transform 1 0 17020 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_180
timestamp 1644511149
transform 1 0 17664 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_205
timestamp 1644511149
transform 1 0 19964 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_212
timestamp 1644511149
transform 1 0 20608 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_219
timestamp 1644511149
transform 1 0 21252 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1644511149
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_274
timestamp 1644511149
transform 1 0 26312 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_81_284
timestamp 1644511149
transform 1 0 27232 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_313
timestamp 1644511149
transform 1 0 29900 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_320
timestamp 1644511149
transform 1 0 30544 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_327
timestamp 1644511149
transform 1 0 31188 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_341
timestamp 1644511149
transform 1 0 32476 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_363
timestamp 1644511149
transform 1 0 34500 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_388
timestamp 1644511149
transform 1 0 36800 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_398
timestamp 1644511149
transform 1 0 37720 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_406
timestamp 1644511149
transform 1 0 38456 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_24
timestamp 1644511149
transform 1 0 3312 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_29
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_52
timestamp 1644511149
transform 1 0 5888 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_57
timestamp 1644511149
transform 1 0 6348 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_80
timestamp 1644511149
transform 1 0 8464 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_88
timestamp 1644511149
transform 1 0 9200 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_95
timestamp 1644511149
transform 1 0 9844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_107
timestamp 1644511149
transform 1 0 10948 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_111
timestamp 1644511149
transform 1 0 11316 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_113
timestamp 1644511149
transform 1 0 11500 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_125
timestamp 1644511149
transform 1 0 12604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_137
timestamp 1644511149
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_169
timestamp 1644511149
transform 1 0 16652 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_192
timestamp 1644511149
transform 1 0 18768 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_205
timestamp 1644511149
transform 1 0 19964 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_82_211
timestamp 1644511149
transform 1 0 20516 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_218
timestamp 1644511149
transform 1 0 21160 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_225
timestamp 1644511149
transform 1 0 21804 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_82_232
timestamp 1644511149
transform 1 0 22448 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_244
timestamp 1644511149
transform 1 0 23552 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_256
timestamp 1644511149
transform 1 0 24656 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_268
timestamp 1644511149
transform 1 0 25760 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_281
timestamp 1644511149
transform 1 0 26956 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_82_289
timestamp 1644511149
transform 1 0 27692 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_295
timestamp 1644511149
transform 1 0 28244 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1644511149
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_330
timestamp 1644511149
transform 1 0 31464 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_82_358
timestamp 1644511149
transform 1 0 34040 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_380
timestamp 1644511149
transform 1 0 36064 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_387
timestamp 1644511149
transform 1 0 36708 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_391
timestamp 1644511149
transform 1 0 37076 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_82_393
timestamp 1644511149
transform 1 0 37260 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_82_399
timestamp 1644511149
transform 1 0 37812 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 38824 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 38824 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 38824 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 38824 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 38824 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 38824 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 38824 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 38824 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 38824 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 38824 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 38824 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 38824 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 38824 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 38824 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 38824 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 38824 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 38824 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 38824 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0708_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12880 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0709_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15088 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  _0710_
timestamp 1644511149
transform 1 0 31832 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0711_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1644511149
transform -1 0 2208 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1644511149
transform -1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0714_
timestamp 1644511149
transform -1 0 2392 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1644511149
transform 1 0 32660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0716_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0718_
timestamp 1644511149
transform 1 0 37352 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0719_
timestamp 1644511149
transform -1 0 2668 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0720_
timestamp 1644511149
transform 1 0 37352 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0722_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8280 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  _0723_
timestamp 1644511149
transform 1 0 9660 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0724_
timestamp 1644511149
transform -1 0 2760 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1644511149
transform 1 0 18124 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0726_
timestamp 1644511149
transform 1 0 37352 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0727_
timestamp 1644511149
transform -1 0 2944 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1644511149
transform 1 0 37352 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0729_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9200 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1644511149
transform 1 0 37904 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0731_
timestamp 1644511149
transform -1 0 2484 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0732_
timestamp 1644511149
transform -1 0 20424 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0734_
timestamp 1644511149
transform -1 0 2576 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0735_
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0736_
timestamp 1644511149
transform 1 0 37352 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1644511149
transform -1 0 22724 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0738_
timestamp 1644511149
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1644511149
transform 1 0 37352 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0740_
timestamp 1644511149
transform -1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0741_
timestamp 1644511149
transform 1 0 9568 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0742_
timestamp 1644511149
transform 1 0 37444 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0744_
timestamp 1644511149
transform 1 0 37444 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1644511149
transform -1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0746_
timestamp 1644511149
transform 1 0 37444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0747_
timestamp 1644511149
transform 1 0 9660 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0748_
timestamp 1644511149
transform -1 0 2944 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0749_
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1644511149
transform 1 0 37444 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0751_
timestamp 1644511149
transform 1 0 37352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1644511149
transform -1 0 15364 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0753_
timestamp 1644511149
transform 1 0 14168 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0754_
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0755_
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0756_
timestamp 1644511149
transform -1 0 2300 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1644511149
transform 1 0 15548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0758_
timestamp 1644511149
transform -1 0 2300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0759_
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0760_
timestamp 1644511149
transform 1 0 14812 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1644511149
transform -1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1644511149
transform -1 0 2208 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0763_
timestamp 1644511149
transform 1 0 35604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0764_
timestamp 1644511149
transform 1 0 35696 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1644511149
transform -1 0 2208 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0766_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 14444 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0767_
timestamp 1644511149
transform 1 0 31372 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1644511149
transform 1 0 31004 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0769_
timestamp 1644511149
transform 1 0 14260 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1644511149
transform -1 0 2944 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1644511149
transform 1 0 30820 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0772_
timestamp 1644511149
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1644511149
transform -1 0 28244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0774_
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0775_
timestamp 1644511149
transform 1 0 23644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1644511149
transform -1 0 28796 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0777_
timestamp 1644511149
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0778_
timestamp 1644511149
transform 1 0 15272 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0779_
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0780_
timestamp 1644511149
transform -1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1644511149
transform 1 0 37444 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1644511149
transform 1 0 37444 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0783_
timestamp 1644511149
transform 1 0 37444 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0784_
timestamp 1644511149
transform -1 0 8096 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0785_
timestamp 1644511149
transform 1 0 7912 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0786_
timestamp 1644511149
transform 1 0 8832 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1644511149
transform 1 0 37352 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1644511149
transform 1 0 37352 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1644511149
transform -1 0 3036 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0790_
timestamp 1644511149
transform -1 0 35236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0791_
timestamp 1644511149
transform 1 0 7912 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0792_
timestamp 1644511149
transform -1 0 2300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0794_
timestamp 1644511149
transform 1 0 22172 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0795_
timestamp 1644511149
transform 1 0 32660 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1644511149
transform -1 0 2392 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0797_
timestamp 1644511149
transform 1 0 7912 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1644511149
transform 1 0 9752 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0799_
timestamp 1644511149
transform 1 0 5612 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1644511149
transform -1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1644511149
transform -1 0 9476 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0802_
timestamp 1644511149
transform 1 0 6532 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0803_
timestamp 1644511149
transform 1 0 7636 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1644511149
transform -1 0 7452 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0805_
timestamp 1644511149
transform 1 0 37444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1644511149
transform 1 0 37444 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0807_
timestamp 1644511149
transform 1 0 11684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1644511149
transform 1 0 37444 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0809_
timestamp 1644511149
transform 1 0 7912 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1644511149
transform 1 0 26220 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0811_
timestamp 1644511149
transform 1 0 37352 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1644511149
transform 1 0 8096 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0813_
timestamp 1644511149
transform 1 0 37352 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1644511149
transform -1 0 7544 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0815_
timestamp 1644511149
transform -1 0 15732 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1644511149
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0817_
timestamp 1644511149
transform -1 0 17480 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0818_
timestamp 1644511149
transform -1 0 19504 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1644511149
transform 1 0 37352 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1644511149
transform 1 0 37352 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0821_
timestamp 1644511149
transform -1 0 15548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1644511149
transform -1 0 2484 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1644511149
transform -1 0 36432 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0825_
timestamp 1644511149
transform -1 0 4048 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0826_
timestamp 1644511149
transform -1 0 4784 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0827_
timestamp 1644511149
transform 1 0 16100 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0828_
timestamp 1644511149
transform 1 0 37904 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1644511149
transform -1 0 2116 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0830_
timestamp 1644511149
transform -1 0 37536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1644511149
transform -1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0832_
timestamp 1644511149
transform -1 0 2208 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0833_
timestamp 1644511149
transform 1 0 13616 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0834_
timestamp 1644511149
transform 1 0 36432 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0835_
timestamp 1644511149
transform -1 0 1656 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0836_
timestamp 1644511149
transform -1 0 35788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0837_
timestamp 1644511149
transform -1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0838_
timestamp 1644511149
transform 1 0 1840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1644511149
transform -1 0 20608 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0840_
timestamp 1644511149
transform 1 0 23000 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1644511149
transform 1 0 33212 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1644511149
transform 1 0 29624 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0843_
timestamp 1644511149
transform 1 0 29624 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1644511149
transform 1 0 28612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1644511149
transform 1 0 28336 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0846_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 36432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0847_
timestamp 1644511149
transform -1 0 37996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1644511149
transform 1 0 28520 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0849_
timestamp 1644511149
transform 1 0 28520 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0850_
timestamp 1644511149
transform -1 0 33120 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0851_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0852_
timestamp 1644511149
transform 1 0 30268 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1644511149
transform -1 0 30912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0854_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29624 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 30268 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1644511149
transform 1 0 28152 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 29072 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0859_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28612 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _0860_
timestamp 1644511149
transform 1 0 29440 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0861_
timestamp 1644511149
transform -1 0 30268 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _0862_
timestamp 1644511149
transform 1 0 29900 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0863_
timestamp 1644511149
transform 1 0 30268 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1644511149
transform -1 0 32200 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0865_
timestamp 1644511149
transform -1 0 32660 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0866_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32476 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _0867_
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0868_
timestamp 1644511149
transform 1 0 31096 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0869_
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1644511149
transform -1 0 16192 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1644511149
transform -1 0 19504 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1644511149
transform -1 0 19504 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1644511149
transform -1 0 21712 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0874_
timestamp 1644511149
transform -1 0 20424 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1644511149
transform 1 0 22080 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0876_
timestamp 1644511149
transform 1 0 22540 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1644511149
transform -1 0 23184 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1644511149
transform -1 0 23460 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0879_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22172 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0880_
timestamp 1644511149
transform -1 0 22632 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0881_
timestamp 1644511149
transform -1 0 21344 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _0882_
timestamp 1644511149
transform -1 0 20148 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0883_
timestamp 1644511149
transform -1 0 19136 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0884_
timestamp 1644511149
transform -1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0885_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16100 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0886_
timestamp 1644511149
transform 1 0 28428 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _0887_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15640 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0888_
timestamp 1644511149
transform 1 0 30176 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _0889_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31280 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform -1 0 30820 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform -1 0 30544 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 28796 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform -1 0 27692 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0894_
timestamp 1644511149
transform 1 0 26864 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0895_
timestamp 1644511149
transform 1 0 27048 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0896_
timestamp 1644511149
transform -1 0 25576 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 25944 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0898_
timestamp 1644511149
transform -1 0 25024 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _0899_
timestamp 1644511149
transform -1 0 25484 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0900_
timestamp 1644511149
transform -1 0 23828 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0901_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25116 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0902_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24564 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0903_
timestamp 1644511149
transform -1 0 26496 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0904_
timestamp 1644511149
transform -1 0 24932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0905_
timestamp 1644511149
transform 1 0 25300 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0906_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25852 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0907_
timestamp 1644511149
transform -1 0 29900 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _0908_
timestamp 1644511149
transform 1 0 27968 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 1644511149
transform -1 0 28612 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0910_
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _0911_
timestamp 1644511149
transform 1 0 29440 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0912_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30268 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0913_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 31188 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0914_
timestamp 1644511149
transform -1 0 28428 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0915_
timestamp 1644511149
transform 1 0 24748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0916_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 24840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0917_
timestamp 1644511149
transform -1 0 28152 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0918_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28152 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0919_
timestamp 1644511149
transform 1 0 26588 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0920_
timestamp 1644511149
transform -1 0 27508 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26036 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0922_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0923_
timestamp 1644511149
transform -1 0 31648 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0924_
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0925_
timestamp 1644511149
transform 1 0 23000 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0926_
timestamp 1644511149
transform 1 0 26496 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0927_
timestamp 1644511149
transform 1 0 27784 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0928_
timestamp 1644511149
transform -1 0 27600 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0929_
timestamp 1644511149
transform 1 0 26404 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0930_
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0931_
timestamp 1644511149
transform -1 0 27416 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0932_
timestamp 1644511149
transform -1 0 26496 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0933_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0934_
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0935_
timestamp 1644511149
transform -1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0936_
timestamp 1644511149
transform 1 0 28060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0937_
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0938_
timestamp 1644511149
transform 1 0 28520 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0939_
timestamp 1644511149
transform 1 0 23000 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0940_
timestamp 1644511149
transform 1 0 23552 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0941_
timestamp 1644511149
transform 1 0 23000 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0942_
timestamp 1644511149
transform 1 0 22080 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0943_
timestamp 1644511149
transform 1 0 23552 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0944_
timestamp 1644511149
transform -1 0 23184 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0945_
timestamp 1644511149
transform 1 0 21804 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0946_
timestamp 1644511149
transform -1 0 20332 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0947_
timestamp 1644511149
transform -1 0 18676 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0948_
timestamp 1644511149
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0949_
timestamp 1644511149
transform -1 0 20976 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0950_
timestamp 1644511149
transform -1 0 19964 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0951_
timestamp 1644511149
transform -1 0 19688 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0952_
timestamp 1644511149
transform -1 0 19504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0953_
timestamp 1644511149
transform 1 0 17204 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0954_
timestamp 1644511149
transform 1 0 18400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0955_
timestamp 1644511149
transform 1 0 17480 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0956_
timestamp 1644511149
transform -1 0 18308 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0957_
timestamp 1644511149
transform 1 0 17480 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0958_
timestamp 1644511149
transform -1 0 16928 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0959_
timestamp 1644511149
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0960_
timestamp 1644511149
transform 1 0 15272 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0961_
timestamp 1644511149
transform 1 0 25024 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _0962_
timestamp 1644511149
transform -1 0 24656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _0963_
timestamp 1644511149
transform 1 0 30268 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0964_
timestamp 1644511149
transform -1 0 26220 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0965_
timestamp 1644511149
transform 1 0 24932 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _0966_
timestamp 1644511149
transform 1 0 31280 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0967_
timestamp 1644511149
transform -1 0 25208 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0968_
timestamp 1644511149
transform -1 0 25668 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0969_
timestamp 1644511149
transform -1 0 24840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0970_
timestamp 1644511149
transform 1 0 26772 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0971_
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0972_
timestamp 1644511149
transform 1 0 27600 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0973_
timestamp 1644511149
transform 1 0 27324 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0974_
timestamp 1644511149
transform 1 0 27140 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0975_
timestamp 1644511149
transform -1 0 28520 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0976_
timestamp 1644511149
transform 1 0 28336 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0977_
timestamp 1644511149
transform 1 0 28888 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0978_
timestamp 1644511149
transform 1 0 29256 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0979_
timestamp 1644511149
transform -1 0 29072 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0980_
timestamp 1644511149
transform 1 0 29440 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0981_
timestamp 1644511149
transform 1 0 31372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0982_
timestamp 1644511149
transform 1 0 30452 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0983_
timestamp 1644511149
transform 1 0 32016 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0984_
timestamp 1644511149
transform -1 0 33120 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0985_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32568 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _0986_
timestamp 1644511149
transform 1 0 33120 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0987_
timestamp 1644511149
transform -1 0 35144 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0988_
timestamp 1644511149
transform -1 0 34684 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0989_
timestamp 1644511149
transform -1 0 34132 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _0990_
timestamp 1644511149
transform -1 0 33764 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0991_
timestamp 1644511149
transform 1 0 32476 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0992_
timestamp 1644511149
transform 1 0 30544 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0993_
timestamp 1644511149
transform 1 0 31004 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0994_
timestamp 1644511149
transform 1 0 33488 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _0995_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33488 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0996_
timestamp 1644511149
transform -1 0 35236 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _0997_
timestamp 1644511149
transform -1 0 35604 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _0998_
timestamp 1644511149
transform 1 0 33488 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0999_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1000_
timestamp 1644511149
transform -1 0 34040 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1001_
timestamp 1644511149
transform -1 0 32292 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1002_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1003_
timestamp 1644511149
transform 1 0 33120 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1004_
timestamp 1644511149
transform 1 0 20976 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1005_
timestamp 1644511149
transform 1 0 23092 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1006_
timestamp 1644511149
transform 1 0 31372 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1007_
timestamp 1644511149
transform 1 0 33304 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1008_
timestamp 1644511149
transform -1 0 33120 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 36432 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1644511149
transform -1 0 34776 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1011_
timestamp 1644511149
transform -1 0 35420 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1012_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35420 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1013_
timestamp 1644511149
transform -1 0 34224 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1014_
timestamp 1644511149
transform -1 0 34408 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1015_
timestamp 1644511149
transform -1 0 36156 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1016_
timestamp 1644511149
transform -1 0 35052 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1017_
timestamp 1644511149
transform 1 0 33672 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1018_
timestamp 1644511149
transform -1 0 33304 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1019_
timestamp 1644511149
transform 1 0 33396 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1020_
timestamp 1644511149
transform 1 0 35236 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1021_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1022_
timestamp 1644511149
transform -1 0 35880 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1023_
timestamp 1644511149
transform 1 0 33764 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1024_
timestamp 1644511149
transform 1 0 34408 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1025_
timestamp 1644511149
transform 1 0 33856 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1026_
timestamp 1644511149
transform -1 0 35696 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1027_
timestamp 1644511149
transform -1 0 34684 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1028_
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1029_
timestamp 1644511149
transform -1 0 35328 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1030_
timestamp 1644511149
transform -1 0 33120 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1031_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 33396 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1032_
timestamp 1644511149
transform -1 0 32476 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1033_
timestamp 1644511149
transform 1 0 32660 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1034_
timestamp 1644511149
transform 1 0 33120 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1035_
timestamp 1644511149
transform 1 0 34224 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1036_
timestamp 1644511149
transform 1 0 33580 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1037_
timestamp 1644511149
transform -1 0 32752 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1038_
timestamp 1644511149
transform 1 0 32108 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1039_
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1040_
timestamp 1644511149
transform 1 0 32292 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1041_
timestamp 1644511149
transform 1 0 30728 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1042_
timestamp 1644511149
transform -1 0 32108 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1043_
timestamp 1644511149
transform -1 0 31096 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1044_
timestamp 1644511149
transform -1 0 31648 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1045_
timestamp 1644511149
transform -1 0 20700 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1046_
timestamp 1644511149
transform 1 0 19320 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1047_
timestamp 1644511149
transform 1 0 32936 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1048_
timestamp 1644511149
transform -1 0 34040 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1049_
timestamp 1644511149
transform -1 0 21252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1050_
timestamp 1644511149
transform 1 0 20608 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1051_
timestamp 1644511149
transform 1 0 19872 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1052_
timestamp 1644511149
transform -1 0 21896 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1053_
timestamp 1644511149
transform 1 0 20608 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1054_
timestamp 1644511149
transform 1 0 20148 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1055_
timestamp 1644511149
transform -1 0 18032 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1056_
timestamp 1644511149
transform 1 0 19136 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1057_
timestamp 1644511149
transform -1 0 23276 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1058_
timestamp 1644511149
transform 1 0 22724 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _1059_
timestamp 1644511149
transform 1 0 20516 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1060_
timestamp 1644511149
transform 1 0 21620 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1061_
timestamp 1644511149
transform -1 0 20056 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1062_
timestamp 1644511149
transform 1 0 16468 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1063_
timestamp 1644511149
transform -1 0 20976 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1064_
timestamp 1644511149
transform 1 0 20516 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1065_
timestamp 1644511149
transform -1 0 22080 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1066_
timestamp 1644511149
transform 1 0 21712 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1067_
timestamp 1644511149
transform 1 0 22632 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1068_
timestamp 1644511149
transform 1 0 22632 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1069_
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1070_
timestamp 1644511149
transform -1 0 22356 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1071_
timestamp 1644511149
transform 1 0 20424 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1072_
timestamp 1644511149
transform -1 0 21988 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1073_
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1074_
timestamp 1644511149
transform 1 0 20424 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1075_
timestamp 1644511149
transform 1 0 21436 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1076_
timestamp 1644511149
transform 1 0 20148 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1077_
timestamp 1644511149
transform 1 0 20884 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1078_
timestamp 1644511149
transform 1 0 20148 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1079_
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1080_
timestamp 1644511149
transform 1 0 20792 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1081_
timestamp 1644511149
transform -1 0 20516 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1082_
timestamp 1644511149
transform 1 0 21896 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1083_
timestamp 1644511149
transform 1 0 20884 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1084_
timestamp 1644511149
transform 1 0 20516 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1085_
timestamp 1644511149
transform 1 0 18032 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1086_
timestamp 1644511149
transform 1 0 18308 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1087_
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1088_
timestamp 1644511149
transform -1 0 19228 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1089_
timestamp 1644511149
transform 1 0 18032 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1090_
timestamp 1644511149
transform 1 0 17112 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1091_
timestamp 1644511149
transform -1 0 19964 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1092_
timestamp 1644511149
transform 1 0 18032 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1093_
timestamp 1644511149
transform 1 0 19228 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1094_
timestamp 1644511149
transform 1 0 18308 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1095_
timestamp 1644511149
transform 1 0 15824 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1096_
timestamp 1644511149
transform 1 0 19044 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1097_
timestamp 1644511149
transform 1 0 18032 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1098_
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1099_
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1100_
timestamp 1644511149
transform 1 0 17296 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1101_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1102_
timestamp 1644511149
transform 1 0 16836 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1103_
timestamp 1644511149
transform 1 0 15272 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1104_
timestamp 1644511149
transform 1 0 15640 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1105_
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1106_
timestamp 1644511149
transform 1 0 16284 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a311oi_1  _1107_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 16100 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1108_
timestamp 1644511149
transform -1 0 23920 0 1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1109_
timestamp 1644511149
transform 1 0 22724 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1110_
timestamp 1644511149
transform -1 0 21252 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1111_
timestamp 1644511149
transform -1 0 20884 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1112_
timestamp 1644511149
transform -1 0 25208 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1113_
timestamp 1644511149
transform -1 0 26128 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1114_
timestamp 1644511149
transform -1 0 25208 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1115_
timestamp 1644511149
transform -1 0 25852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1116_
timestamp 1644511149
transform -1 0 25392 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1644511149
transform -1 0 25484 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1118_
timestamp 1644511149
transform 1 0 25208 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1119_
timestamp 1644511149
transform 1 0 25944 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1120_
timestamp 1644511149
transform 1 0 23920 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1121_
timestamp 1644511149
transform -1 0 23276 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1122_
timestamp 1644511149
transform -1 0 29808 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and4b_1  _1123_
timestamp 1644511149
transform 1 0 24472 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1124_
timestamp 1644511149
transform -1 0 26312 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1125_
timestamp 1644511149
transform 1 0 25760 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1126_
timestamp 1644511149
transform 1 0 27324 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1127_
timestamp 1644511149
transform -1 0 24656 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1128_
timestamp 1644511149
transform -1 0 25392 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1129_
timestamp 1644511149
transform -1 0 23368 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1644511149
transform -1 0 23920 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1131_
timestamp 1644511149
transform 1 0 23552 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1132_
timestamp 1644511149
transform 1 0 22632 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1133_
timestamp 1644511149
transform -1 0 23092 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1134_
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1135_
timestamp 1644511149
transform 1 0 23736 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1136_
timestamp 1644511149
transform 1 0 22356 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1137_
timestamp 1644511149
transform 1 0 23092 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1138_
timestamp 1644511149
transform 1 0 23460 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1139_
timestamp 1644511149
transform 1 0 23368 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1140_
timestamp 1644511149
transform -1 0 23092 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1141_
timestamp 1644511149
transform -1 0 25760 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1142_
timestamp 1644511149
transform -1 0 25208 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1143_
timestamp 1644511149
transform -1 0 24748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1144_
timestamp 1644511149
transform 1 0 24472 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1145_
timestamp 1644511149
transform 1 0 30360 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1146_
timestamp 1644511149
transform 1 0 24472 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1147_
timestamp 1644511149
transform -1 0 24932 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1148_
timestamp 1644511149
transform -1 0 26220 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1149_
timestamp 1644511149
transform -1 0 27324 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1150_
timestamp 1644511149
transform -1 0 27600 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1151_
timestamp 1644511149
transform -1 0 26496 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1152_
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1153_
timestamp 1644511149
transform -1 0 27416 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1154_
timestamp 1644511149
transform 1 0 28980 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1155_
timestamp 1644511149
transform 1 0 27876 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1156_
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1157_
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1158_
timestamp 1644511149
transform -1 0 21988 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1159_
timestamp 1644511149
transform 1 0 29900 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1160_
timestamp 1644511149
transform 1 0 30544 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1161_
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1162_
timestamp 1644511149
transform -1 0 27416 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1163_
timestamp 1644511149
transform -1 0 26312 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1164_
timestamp 1644511149
transform 1 0 27876 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1165_
timestamp 1644511149
transform 1 0 27692 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1166_
timestamp 1644511149
transform 1 0 26680 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1167_
timestamp 1644511149
transform 1 0 26036 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1168_
timestamp 1644511149
transform -1 0 27692 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1169_
timestamp 1644511149
transform -1 0 27600 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1170_
timestamp 1644511149
transform 1 0 28428 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1171_
timestamp 1644511149
transform 1 0 28704 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1172_
timestamp 1644511149
transform 1 0 29716 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1173_
timestamp 1644511149
transform -1 0 30084 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1174_
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1175_
timestamp 1644511149
transform -1 0 28612 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1176_
timestamp 1644511149
transform 1 0 30728 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1177_
timestamp 1644511149
transform 1 0 31372 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1178_
timestamp 1644511149
transform -1 0 32108 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1179_
timestamp 1644511149
transform -1 0 31648 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1180_
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1181_
timestamp 1644511149
transform -1 0 33120 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1182_
timestamp 1644511149
transform 1 0 32016 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1183_
timestamp 1644511149
transform 1 0 32660 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1184_
timestamp 1644511149
transform 1 0 33948 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1185_
timestamp 1644511149
transform -1 0 34684 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1186_
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1187_
timestamp 1644511149
transform -1 0 36248 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1188_
timestamp 1644511149
transform -1 0 34224 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1189_
timestamp 1644511149
transform 1 0 35052 0 -1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1190_
timestamp 1644511149
transform 1 0 35604 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1191_
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1192_
timestamp 1644511149
transform -1 0 27232 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1193_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35328 0 1 39168
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1194_
timestamp 1644511149
transform 1 0 32292 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1195_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32292 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1196_
timestamp 1644511149
transform -1 0 35236 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1197_
timestamp 1644511149
transform -1 0 33672 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 32568 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1199_
timestamp 1644511149
transform 1 0 35420 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1200_
timestamp 1644511149
transform 1 0 35604 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1201_
timestamp 1644511149
transform -1 0 35144 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1202_
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1203_
timestamp 1644511149
transform -1 0 34316 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1204_
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1205_
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1206_
timestamp 1644511149
transform -1 0 35144 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1207_
timestamp 1644511149
transform -1 0 34960 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1208_
timestamp 1644511149
transform -1 0 36984 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1209_
timestamp 1644511149
transform -1 0 36248 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1210_
timestamp 1644511149
transform 1 0 37352 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1211_
timestamp 1644511149
transform 1 0 37352 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1212_
timestamp 1644511149
transform -1 0 36340 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1213_
timestamp 1644511149
transform -1 0 35512 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1214_
timestamp 1644511149
transform -1 0 37720 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1215_
timestamp 1644511149
transform 1 0 36432 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1216_
timestamp 1644511149
transform -1 0 36340 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1217_
timestamp 1644511149
transform -1 0 36616 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1218_
timestamp 1644511149
transform -1 0 35788 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1219_
timestamp 1644511149
transform -1 0 37812 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1220_
timestamp 1644511149
transform 1 0 34224 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _1221_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 33488 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1222_
timestamp 1644511149
transform -1 0 14536 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1223_
timestamp 1644511149
transform -1 0 14352 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1224_
timestamp 1644511149
transform 1 0 17296 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1225_
timestamp 1644511149
transform -1 0 15824 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1226_
timestamp 1644511149
transform -1 0 14536 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1227_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1228_
timestamp 1644511149
transform -1 0 17756 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1229_
timestamp 1644511149
transform -1 0 15824 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1230_
timestamp 1644511149
transform 1 0 14720 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1231_
timestamp 1644511149
transform -1 0 15824 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1232_
timestamp 1644511149
transform 1 0 15180 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1233_
timestamp 1644511149
transform -1 0 17112 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1234_
timestamp 1644511149
transform 1 0 15916 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1235_
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1236_
timestamp 1644511149
transform -1 0 17848 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1237_
timestamp 1644511149
transform 1 0 17204 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1238_
timestamp 1644511149
transform 1 0 18216 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1239_
timestamp 1644511149
transform -1 0 19504 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1240_
timestamp 1644511149
transform 1 0 17848 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1241_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1242_
timestamp 1644511149
transform 1 0 16468 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1243_
timestamp 1644511149
transform -1 0 18308 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1244_
timestamp 1644511149
transform 1 0 17940 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1245_
timestamp 1644511149
transform 1 0 18032 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1246_
timestamp 1644511149
transform -1 0 17296 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1247_
timestamp 1644511149
transform -1 0 16468 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1248_
timestamp 1644511149
transform -1 0 17204 0 1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1249_
timestamp 1644511149
transform -1 0 16744 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1250_
timestamp 1644511149
transform -1 0 17112 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1251_
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1252_
timestamp 1644511149
transform -1 0 18952 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1253_
timestamp 1644511149
transform 1 0 16744 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1254_
timestamp 1644511149
transform -1 0 19780 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1255_
timestamp 1644511149
transform -1 0 18768 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1256_
timestamp 1644511149
transform -1 0 18216 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1257_
timestamp 1644511149
transform 1 0 20332 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1258_
timestamp 1644511149
transform -1 0 21068 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1259_
timestamp 1644511149
transform 1 0 20792 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1260_
timestamp 1644511149
transform -1 0 21344 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1261_
timestamp 1644511149
transform -1 0 19688 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1262_
timestamp 1644511149
transform 1 0 19320 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1263_
timestamp 1644511149
transform 1 0 20056 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1264_
timestamp 1644511149
transform 1 0 17480 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1265_
timestamp 1644511149
transform 1 0 17572 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1266_
timestamp 1644511149
transform -1 0 20424 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1267_
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1268_
timestamp 1644511149
transform 1 0 20424 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1269_
timestamp 1644511149
transform 1 0 16376 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1270_
timestamp 1644511149
transform 1 0 17204 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1271_
timestamp 1644511149
transform 1 0 18216 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1272_
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1273_
timestamp 1644511149
transform 1 0 21160 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1274_
timestamp 1644511149
transform 1 0 19872 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1275_
timestamp 1644511149
transform -1 0 20976 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1276_
timestamp 1644511149
transform 1 0 19044 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1277_
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1278_
timestamp 1644511149
transform 1 0 19504 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1279_
timestamp 1644511149
transform -1 0 20240 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1280_
timestamp 1644511149
transform 1 0 20792 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1281_
timestamp 1644511149
transform 1 0 20976 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1282_
timestamp 1644511149
transform 1 0 21620 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1283_
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1284_
timestamp 1644511149
transform 1 0 22632 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1285_
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1286_
timestamp 1644511149
transform 1 0 25300 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1287_
timestamp 1644511149
transform 1 0 22632 0 1 44608
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1288_
timestamp 1644511149
transform 1 0 19964 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1289_
timestamp 1644511149
transform 1 0 19872 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1290_
timestamp 1644511149
transform -1 0 22724 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1291_
timestamp 1644511149
transform 1 0 22448 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1292_
timestamp 1644511149
transform 1 0 22080 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1293_
timestamp 1644511149
transform 1 0 23460 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1294_
timestamp 1644511149
transform -1 0 24012 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1295_
timestamp 1644511149
transform -1 0 26220 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1296_
timestamp 1644511149
transform 1 0 25116 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1297_
timestamp 1644511149
transform -1 0 26312 0 -1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1298_
timestamp 1644511149
transform 1 0 25760 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1299_
timestamp 1644511149
transform -1 0 27600 0 1 44608
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1300_
timestamp 1644511149
transform -1 0 27232 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1301_
timestamp 1644511149
transform 1 0 26772 0 1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1302_
timestamp 1644511149
transform -1 0 28060 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1303_
timestamp 1644511149
transform 1 0 29532 0 -1 43520
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1304_
timestamp 1644511149
transform 1 0 29716 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1305_
timestamp 1644511149
transform 1 0 30360 0 -1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1306_
timestamp 1644511149
transform -1 0 31372 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1307_
timestamp 1644511149
transform -1 0 29992 0 1 41344
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1308_
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1309_
timestamp 1644511149
transform -1 0 30176 0 1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1310_
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1311_
timestamp 1644511149
transform 1 0 26772 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1312_
timestamp 1644511149
transform -1 0 29900 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1313_
timestamp 1644511149
transform -1 0 28152 0 1 42432
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _1314_
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  _1315_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1316_
timestamp 1644511149
transform -1 0 28796 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1317_
timestamp 1644511149
transform 1 0 25024 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1318_
timestamp 1644511149
transform 1 0 25024 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1319_
timestamp 1644511149
transform 1 0 25024 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1320_
timestamp 1644511149
transform 1 0 25760 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1321_
timestamp 1644511149
transform 1 0 27968 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1322_
timestamp 1644511149
transform 1 0 28428 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1323_
timestamp 1644511149
transform -1 0 24564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1324_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1325_
timestamp 1644511149
transform -1 0 25116 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1326_
timestamp 1644511149
transform -1 0 21344 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1327_
timestamp 1644511149
transform -1 0 19504 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1328_
timestamp 1644511149
transform 1 0 17020 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1329_
timestamp 1644511149
transform 1 0 16008 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1330_
timestamp 1644511149
transform 1 0 14168 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1331_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1332_
timestamp 1644511149
transform 1 0 24656 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1333_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1334_
timestamp 1644511149
transform -1 0 28428 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1335_
timestamp 1644511149
transform 1 0 26680 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1336_
timestamp 1644511149
transform -1 0 29900 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1337_
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1338_
timestamp 1644511149
transform 1 0 30176 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1339_
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1340_
timestamp 1644511149
transform -1 0 30636 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1341_
timestamp 1644511149
transform 1 0 31280 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1342_
timestamp 1644511149
transform 1 0 34868 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1343_
timestamp 1644511149
transform 1 0 35236 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1344_
timestamp 1644511149
transform 1 0 35052 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1345_
timestamp 1644511149
transform 1 0 32936 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1346_
timestamp 1644511149
transform -1 0 32660 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1347_
timestamp 1644511149
transform -1 0 31648 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1348_
timestamp 1644511149
transform 1 0 18400 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1349_
timestamp 1644511149
transform 1 0 34040 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1350_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22356 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _1351_
timestamp 1644511149
transform 1 0 22448 0 -1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1352_
timestamp 1644511149
transform 1 0 19872 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1353_
timestamp 1644511149
transform -1 0 23828 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1354_
timestamp 1644511149
transform 1 0 17940 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1355_
timestamp 1644511149
transform 1 0 17848 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1356_
timestamp 1644511149
transform -1 0 17388 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1357_
timestamp 1644511149
transform 1 0 14444 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1358_
timestamp 1644511149
transform 1 0 22632 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1359_
timestamp 1644511149
transform -1 0 21436 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1360_
timestamp 1644511149
transform 1 0 22080 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1361_
timestamp 1644511149
transform 1 0 22264 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1362_
timestamp 1644511149
transform 1 0 22724 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1363_
timestamp 1644511149
transform 1 0 25024 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1364_
timestamp 1644511149
transform -1 0 28888 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1365_
timestamp 1644511149
transform -1 0 31464 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1366_
timestamp 1644511149
transform 1 0 27416 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1367_
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1368_
timestamp 1644511149
transform 1 0 28796 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1369_
timestamp 1644511149
transform 1 0 30176 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1370_
timestamp 1644511149
transform -1 0 33580 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1371_
timestamp 1644511149
transform -1 0 33580 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1372_
timestamp 1644511149
transform 1 0 32384 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1373_
timestamp 1644511149
transform 1 0 33580 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1374_
timestamp 1644511149
transform 1 0 33948 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1375_
timestamp 1644511149
transform 1 0 35328 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1376_
timestamp 1644511149
transform -1 0 28060 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1377_
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1378_
timestamp 1644511149
transform 1 0 35328 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1379_
timestamp 1644511149
transform 1 0 33948 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1380_
timestamp 1644511149
transform 1 0 32752 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1381_
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1382_
timestamp 1644511149
transform 1 0 36248 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1383_
timestamp 1644511149
transform 1 0 36708 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1384_
timestamp 1644511149
transform 1 0 35328 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1385_
timestamp 1644511149
transform 1 0 36156 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1386_
timestamp 1644511149
transform 1 0 33028 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1387_
timestamp 1644511149
transform 1 0 14352 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1388_
timestamp 1644511149
transform 1 0 14904 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1389_
timestamp 1644511149
transform -1 0 18216 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1390_
timestamp 1644511149
transform 1 0 14260 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1391_
timestamp 1644511149
transform 1 0 14812 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1392_
timestamp 1644511149
transform 1 0 15548 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1393_
timestamp 1644511149
transform 1 0 16928 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1394_
timestamp 1644511149
transform -1 0 20240 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1395_
timestamp 1644511149
transform 1 0 18216 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1396_
timestamp 1644511149
transform 1 0 16192 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1397_
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1398_
timestamp 1644511149
transform 1 0 15456 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1399_
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1400_
timestamp 1644511149
transform 1 0 18492 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1401_
timestamp 1644511149
transform -1 0 21252 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1402_
timestamp 1644511149
transform -1 0 21988 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1403_
timestamp 1644511149
transform 1 0 18584 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1404_
timestamp 1644511149
transform 1 0 19872 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1405_
timestamp 1644511149
transform 1 0 16744 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1406_
timestamp 1644511149
transform 1 0 18032 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1407_
timestamp 1644511149
transform -1 0 21344 0 -1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1408_
timestamp 1644511149
transform 1 0 18124 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1409_
timestamp 1644511149
transform 1 0 19780 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1410_
timestamp 1644511149
transform 1 0 20792 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1411_
timestamp 1644511149
transform -1 0 23644 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1412_
timestamp 1644511149
transform -1 0 24932 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1413_
timestamp 1644511149
transform 1 0 21620 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1414_
timestamp 1644511149
transform 1 0 23920 0 -1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1415_
timestamp 1644511149
transform 1 0 24840 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1416_
timestamp 1644511149
transform 1 0 25300 0 1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1417_
timestamp 1644511149
transform -1 0 28428 0 -1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1418_
timestamp 1644511149
transform 1 0 27600 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1419_
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1420_
timestamp 1644511149
transform -1 0 32292 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1421_
timestamp 1644511149
transform 1 0 28612 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1422_
timestamp 1644511149
transform -1 0 27784 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1423__9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1424__10
timestamp 1644511149
transform -1 0 1840 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1425__11
timestamp 1644511149
transform -1 0 18400 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1426__12
timestamp 1644511149
transform -1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1427__13
timestamp 1644511149
transform -1 0 33580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1428__14
timestamp 1644511149
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1429__15
timestamp 1644511149
transform 1 0 37628 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1430__16
timestamp 1644511149
transform -1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1431__17
timestamp 1644511149
transform 1 0 37904 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1432__18
timestamp 1644511149
transform -1 0 36708 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1433__19
timestamp 1644511149
transform -1 0 36800 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1434__20
timestamp 1644511149
transform 1 0 19320 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1435__21
timestamp 1644511149
transform 1 0 37536 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1436__22
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1437__23
timestamp 1644511149
transform 1 0 17388 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1438__24
timestamp 1644511149
transform 1 0 1840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1439__25
timestamp 1644511149
transform 1 0 37628 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1440__26
timestamp 1644511149
transform -1 0 36800 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1441__27
timestamp 1644511149
transform -1 0 3588 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1442__28
timestamp 1644511149
transform 1 0 37904 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1443__29
timestamp 1644511149
transform 1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1444__30
timestamp 1644511149
transform -1 0 36800 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1445__31
timestamp 1644511149
transform -1 0 22448 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1446__32
timestamp 1644511149
transform -1 0 11040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1447__33
timestamp 1644511149
transform 1 0 37628 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1448__34
timestamp 1644511149
transform 1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1449__35
timestamp 1644511149
transform 1 0 37904 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1450__36
timestamp 1644511149
transform -1 0 1840 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1451__37
timestamp 1644511149
transform 1 0 37628 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1452__38
timestamp 1644511149
transform -1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1453__39
timestamp 1644511149
transform -1 0 36800 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1454__40
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1455__41
timestamp 1644511149
transform -1 0 34132 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1456__42
timestamp 1644511149
transform -1 0 24656 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1457__43
timestamp 1644511149
transform 1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1458__44
timestamp 1644511149
transform -1 0 2116 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1459__45
timestamp 1644511149
transform 1 0 35604 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1460__46
timestamp 1644511149
transform -1 0 15272 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1461__47
timestamp 1644511149
transform -1 0 36800 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1462__48
timestamp 1644511149
transform -1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1463__49
timestamp 1644511149
transform -1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1464__50
timestamp 1644511149
transform -1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1465__51
timestamp 1644511149
transform -1 0 36800 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1466__52
timestamp 1644511149
transform -1 0 1840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1467__53
timestamp 1644511149
transform -1 0 1748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1468__54
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1469__55
timestamp 1644511149
transform -1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1470__56
timestamp 1644511149
transform -1 0 1932 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1471__57
timestamp 1644511149
transform -1 0 31188 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1472__58
timestamp 1644511149
transform 1 0 1932 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1473__59
timestamp 1644511149
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1474__60
timestamp 1644511149
transform 1 0 37904 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1475__61
timestamp 1644511149
transform 1 0 23184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1476__62
timestamp 1644511149
transform -1 0 28244 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1477__63
timestamp 1644511149
transform -1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1478__64
timestamp 1644511149
transform -1 0 29808 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1479__65
timestamp 1644511149
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1480__66
timestamp 1644511149
transform 1 0 37628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1481__67
timestamp 1644511149
transform 1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1482__68
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1483__69
timestamp 1644511149
transform -1 0 2484 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1484__70
timestamp 1644511149
transform 1 0 37628 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1485__71
timestamp 1644511149
transform -1 0 36800 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1486__72
timestamp 1644511149
transform 1 0 35880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1487__73
timestamp 1644511149
transform -1 0 9200 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1488__74
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1489__75
timestamp 1644511149
transform 1 0 22356 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1490__76
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1491__77
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1492__78
timestamp 1644511149
transform 1 0 22172 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1493__79
timestamp 1644511149
transform -1 0 33672 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1494__80
timestamp 1644511149
transform -1 0 2024 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1495__81
timestamp 1644511149
transform -1 0 36800 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1496__82
timestamp 1644511149
transform -1 0 6624 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1497__83
timestamp 1644511149
transform 1 0 4416 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1498__84
timestamp 1644511149
transform -1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1499__85
timestamp 1644511149
transform 1 0 2576 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1500__86
timestamp 1644511149
transform 1 0 37904 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1501__87
timestamp 1644511149
transform -1 0 36800 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1502__88
timestamp 1644511149
transform 1 0 35880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1503__89
timestamp 1644511149
transform -1 0 6624 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1504__90
timestamp 1644511149
transform 1 0 5612 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1505__91
timestamp 1644511149
transform 1 0 37628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1506__92
timestamp 1644511149
transform -1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1507__93
timestamp 1644511149
transform -1 0 27232 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1508__94
timestamp 1644511149
transform 1 0 9568 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1509__95
timestamp 1644511149
transform -1 0 36800 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1510__96
timestamp 1644511149
transform 1 0 7176 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1511__97
timestamp 1644511149
transform 1 0 5060 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1512__98
timestamp 1644511149
transform 1 0 16744 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1513__99
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1514__100
timestamp 1644511149
transform -1 0 37904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1515__101
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1516__102
timestamp 1644511149
transform -1 0 20516 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1517__103
timestamp 1644511149
transform -1 0 36800 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1518__104
timestamp 1644511149
transform 1 0 36524 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1519__105
timestamp 1644511149
transform 1 0 1564 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1520__106
timestamp 1644511149
transform -1 0 38180 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1521__107
timestamp 1644511149
transform 1 0 1564 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1522__108
timestamp 1644511149
transform -1 0 35144 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1523__109
timestamp 1644511149
transform -1 0 5428 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1524__110
timestamp 1644511149
transform -1 0 1840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1525__111
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1526__112
timestamp 1644511149
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1527_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6624 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1528_
timestamp 1644511149
transform 1 0 1564 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1529_
timestamp 1644511149
transform 1 0 18124 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1530_
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1531_
timestamp 1644511149
transform 1 0 33212 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1532_
timestamp 1644511149
transform 1 0 2944 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1533_
timestamp 1644511149
transform -1 0 38180 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1534_
timestamp 1644511149
transform 1 0 1932 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1535_
timestamp 1644511149
transform -1 0 38180 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1536_
timestamp 1644511149
transform 1 0 36248 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1537_
timestamp 1644511149
transform 1 0 36248 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1538_
timestamp 1644511149
transform 1 0 19964 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1539_
timestamp 1644511149
transform -1 0 38180 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1540_
timestamp 1644511149
transform 1 0 2024 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1541_
timestamp 1644511149
transform 1 0 18032 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1542_
timestamp 1644511149
transform 1 0 2024 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1543_
timestamp 1644511149
transform -1 0 38180 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1544_
timestamp 1644511149
transform 1 0 36248 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1545_
timestamp 1644511149
transform -1 0 3312 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1546_
timestamp 1644511149
transform -1 0 38180 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1547_
timestamp 1644511149
transform 1 0 1840 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1548_
timestamp 1644511149
transform 1 0 36248 0 1 43520
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1549_
timestamp 1644511149
transform 1 0 22080 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1550_
timestamp 1644511149
transform 1 0 10396 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1551_
timestamp 1644511149
transform -1 0 38180 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1552_
timestamp 1644511149
transform 1 0 8464 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1553_
timestamp 1644511149
transform -1 0 38180 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1554_
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1555_
timestamp 1644511149
transform -1 0 38180 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1556_
timestamp 1644511149
transform 1 0 4600 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1557_
timestamp 1644511149
transform 1 0 36248 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1558_
timestamp 1644511149
transform -1 0 36800 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1559_
timestamp 1644511149
transform 1 0 32568 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1560_
timestamp 1644511149
transform 1 0 24380 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1561_
timestamp 1644511149
transform 1 0 8924 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1562_
timestamp 1644511149
transform 1 0 1840 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1563_
timestamp 1644511149
transform 1 0 36248 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1564_
timestamp 1644511149
transform 1 0 14904 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1565_
timestamp 1644511149
transform 1 0 36248 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1566_
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1567_
timestamp 1644511149
transform 1 0 16192 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1568_
timestamp 1644511149
transform 1 0 1656 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1569_
timestamp 1644511149
transform 1 0 36248 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1570_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1571_
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1572_
timestamp 1644511149
transform 1 0 35328 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1573_
timestamp 1644511149
transform 1 0 31464 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1574_
timestamp 1644511149
transform -1 0 16192 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1575_
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1576_
timestamp 1644511149
transform 1 0 35604 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1577_
timestamp 1644511149
transform 1 0 34868 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1578_
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1579_
timestamp 1644511149
transform 1 0 30912 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1580_
timestamp 1644511149
transform -1 0 3312 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1581_
timestamp 1644511149
transform 1 0 27784 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1582_
timestamp 1644511149
transform -1 0 38180 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1583_
timestamp 1644511149
transform 1 0 23828 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1584_
timestamp 1644511149
transform 1 0 27968 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1585_
timestamp 1644511149
transform 1 0 2944 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1586_
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1587_
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1588_
timestamp 1644511149
transform -1 0 38180 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1589_
timestamp 1644511149
transform -1 0 3312 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1590_
timestamp 1644511149
transform 1 0 1656 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1591_
timestamp 1644511149
transform 1 0 2024 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1592_
timestamp 1644511149
transform -1 0 38180 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1593_
timestamp 1644511149
transform 1 0 36248 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1594_
timestamp 1644511149
transform 1 0 36248 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1595_
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1596_
timestamp 1644511149
transform -1 0 36800 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1597_
timestamp 1644511149
transform 1 0 23368 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1598_
timestamp 1644511149
transform 1 0 34776 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1599_
timestamp 1644511149
transform 1 0 32108 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1600_
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1601_
timestamp 1644511149
transform 1 0 33396 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1602_
timestamp 1644511149
transform 1 0 1656 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1603_
timestamp 1644511149
transform 1 0 36248 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1604_
timestamp 1644511149
transform 1 0 5796 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1605_
timestamp 1644511149
transform -1 0 5888 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1606_
timestamp 1644511149
transform 1 0 9016 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1607_
timestamp 1644511149
transform -1 0 3312 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1608_
timestamp 1644511149
transform -1 0 38180 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1609_
timestamp 1644511149
transform 1 0 36248 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1610_
timestamp 1644511149
transform 1 0 36248 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1611_
timestamp 1644511149
transform 1 0 6348 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1612_
timestamp 1644511149
transform 1 0 6532 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1613_
timestamp 1644511149
transform -1 0 38180 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1614_
timestamp 1644511149
transform 1 0 11684 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1615_
timestamp 1644511149
transform 1 0 26220 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1616_
timestamp 1644511149
transform -1 0 9844 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1617_
timestamp 1644511149
transform 1 0 36248 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1618_
timestamp 1644511149
transform -1 0 8464 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1619_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1620_
timestamp 1644511149
transform 1 0 16836 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1621_
timestamp 1644511149
transform -1 0 19412 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1622_
timestamp 1644511149
transform -1 0 34224 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1623_
timestamp 1644511149
transform 1 0 36248 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1624_
timestamp 1644511149
transform 1 0 20148 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1625_
timestamp 1644511149
transform 1 0 36248 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1626_
timestamp 1644511149
transform -1 0 36800 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1627_
timestamp 1644511149
transform -1 0 3312 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1628_
timestamp 1644511149
transform -1 0 36800 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1629_
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1630_
timestamp 1644511149
transform -1 0 34224 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1631_
timestamp 1644511149
transform 1 0 3956 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1632_
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1633_
timestamp 1644511149
transform -1 0 3496 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1634_
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform -1 0 27416 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform -1 0 22540 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 20976 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform -1 0 31004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 30544 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform -1 0 20516 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform -1 0 21252 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 31004 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 30636 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input1
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1644511149
transform 1 0 20884 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1644511149
transform 1 0 35880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1644511149
transform -1 0 38180 0 -1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1644511149
transform 1 0 4324 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input8
timestamp 1644511149
transform -1 0 38180 0 -1 13056
box -38 -48 590 592
<< labels >>
rlabel metal3 s 0 41428 800 41668 6 active
port 0 nsew signal input
rlabel metal2 s 13514 0 13626 800 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 19954 49200 20066 50000 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 44828 800 45068 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 39200 42788 40000 43028 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 21242 0 21354 800 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 11582 49200 11694 50000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 39200 44828 40000 45068 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 39200 8788 40000 9028 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 3854 49200 3966 50000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 5786 49200 5898 50000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 38630 0 38742 800 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 0 14228 800 14468 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 0 25788 800 26028 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 16948 800 17188 6 io_in[21]
port 14 nsew signal input
rlabel metal3 s 39200 19668 40000 19908 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 3210 49200 3322 50000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 634 49200 746 50000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 33478 0 33590 800 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 32834 0 32946 800 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 39200 14908 40000 15148 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 29614 0 29726 800 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 39274 49200 39386 50000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 14802 0 14914 800 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 39200 23068 40000 23308 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 40068 800 40308 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 27682 0 27794 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 23068 800 23308 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 28970 49200 29082 50000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 34122 49200 34234 50000 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 39200 33268 40000 33508 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 34766 49200 34878 50000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 20598 49200 20710 50000 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 39200 32588 40000 32828 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 39200 48228 40000 48468 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 0 27828 800 28068 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 0 18988 800 19228 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 39200 35308 40000 35548 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 2566 49200 2678 50000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 23818 0 23930 800 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 0 15588 800 15828 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal3 s 39200 30548 40000 30788 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal3 s 39200 18308 40000 18548 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal3 s 39200 17628 40000 17868 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal3 s 0 4028 800 4268 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal2 s 7074 49200 7186 50000 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 39200 7428 40000 7668 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal2 s 12226 0 12338 800 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal2 s 27038 49200 27150 50000 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal2 s 8362 49200 8474 50000 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal2 s 35410 0 35522 800 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 39200 24428 40000 24668 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal3 s 0 46868 800 47108 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal2 s 4498 0 4610 800 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal2 s 17378 49200 17490 50000 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal2 s 18022 49200 18134 50000 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal3 s 39200 2668 40000 2908 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 39200 40068 40000 40308 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal2 s 21242 49200 21354 50000 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal2 s 37986 0 38098 800 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal3 s 39200 33948 40000 34188 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal2 s 32190 49200 32302 50000 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal3 s 0 47548 800 47788 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal2 s 36698 0 36810 800 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal3 s 0 22388 800 22628 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal3 s 39200 4028 40000 4268 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal2 s 5142 49200 5254 50000 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 0 19668 800 19908 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal3 s 0 10148 800 10388 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 0 16268 800 16508 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal2 s 22530 0 22642 800 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 39200 5388 40000 5628 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 0 29188 800 29428 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal3 s 39200 21028 40000 21268 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal2 s 6430 49200 6542 50000 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal2 s 3854 0 3966 800 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal2 s 9650 0 9762 800 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal3 s 39200 47548 40000 47788 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 39200 29868 40000 30108 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 0 1988 800 2228 6 io_out[11]
port 79 nsew signal tristate
rlabel metal3 s 0 6748 800 6988 6 io_out[12]
port 80 nsew signal tristate
rlabel metal2 s 36054 0 36166 800 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 39200 41428 40000 41668 6 io_out[14]
port 82 nsew signal tristate
rlabel metal3 s 0 37348 800 37588 6 io_out[15]
port 83 nsew signal tristate
rlabel metal3 s 39200 29188 40000 29428 6 io_out[16]
port 84 nsew signal tristate
rlabel metal2 s 36054 49200 36166 50000 6 io_out[17]
port 85 nsew signal tristate
rlabel metal3 s 39200 1988 40000 2228 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 0 21708 800 21948 6 io_out[19]
port 87 nsew signal tristate
rlabel metal2 s 24462 49200 24574 50000 6 io_out[1]
port 88 nsew signal tristate
rlabel metal2 s 31546 49200 31658 50000 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 0 35988 800 36228 6 io_out[21]
port 90 nsew signal tristate
rlabel metal2 s 28326 0 28438 800 6 io_out[22]
port 91 nsew signal tristate
rlabel metal3 s 39200 25788 40000 26028 6 io_out[23]
port 92 nsew signal tristate
rlabel metal2 s 24462 0 24574 800 6 io_out[24]
port 93 nsew signal tristate
rlabel metal2 s 28326 49200 28438 50000 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 0 4708 800 4948 6 io_out[26]
port 95 nsew signal tristate
rlabel metal2 s 29614 49200 29726 50000 6 io_out[27]
port 96 nsew signal tristate
rlabel metal2 s 15446 0 15558 800 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 39200 6068 40000 6308 6 io_out[29]
port 98 nsew signal tristate
rlabel metal2 s 6430 0 6542 800 6 io_out[2]
port 99 nsew signal tristate
rlabel metal3 s 0 5388 800 5628 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 0 12868 800 13108 6 io_out[31]
port 101 nsew signal tristate
rlabel metal3 s 0 42108 800 42348 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 39200 11508 40000 11748 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 39200 42108 40000 42348 6 io_out[34]
port 104 nsew signal tristate
rlabel metal3 s 39200 39388 40000 39628 6 io_out[35]
port 105 nsew signal tristate
rlabel metal2 s 9006 49200 9118 50000 6 io_out[36]
port 106 nsew signal tristate
rlabel metal3 s 39200 45508 40000 45748 6 io_out[37]
port 107 nsew signal tristate
rlabel metal3 s 0 38708 800 38948 6 io_out[3]
port 108 nsew signal tristate
rlabel metal3 s 39200 31908 40000 32148 6 io_out[4]
port 109 nsew signal tristate
rlabel metal2 s 15446 49200 15558 50000 6 io_out[5]
port 110 nsew signal tristate
rlabel metal2 s 37986 49200 38098 50000 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 0 17628 800 17868 6 io_out[7]
port 112 nsew signal tristate
rlabel metal2 s 16734 0 16846 800 6 io_out[8]
port 113 nsew signal tristate
rlabel metal3 s 0 13548 800 13788 6 io_out[9]
port 114 nsew signal tristate
rlabel metal3 s 39200 12188 40000 12428 6 la1_data_in[0]
port 115 nsew signal input
rlabel metal2 s 19310 0 19422 800 6 la1_data_in[10]
port 116 nsew signal input
rlabel metal3 s 39200 10828 40000 11068 6 la1_data_in[11]
port 117 nsew signal input
rlabel metal3 s 0 33948 800 34188 6 la1_data_in[12]
port 118 nsew signal input
rlabel metal2 s 30258 0 30370 800 6 la1_data_in[13]
port 119 nsew signal input
rlabel metal3 s 0 11508 800 11748 6 la1_data_in[14]
port 120 nsew signal input
rlabel metal2 s 9650 49200 9762 50000 6 la1_data_in[15]
port 121 nsew signal input
rlabel metal2 s 23174 49200 23286 50000 6 la1_data_in[16]
port 122 nsew signal input
rlabel metal2 s 16734 49200 16846 50000 6 la1_data_in[17]
port 123 nsew signal input
rlabel metal2 s 39274 0 39386 800 6 la1_data_in[18]
port 124 nsew signal input
rlabel metal2 s 10938 49200 11050 50000 6 la1_data_in[19]
port 125 nsew signal input
rlabel metal2 s 18022 0 18134 800 6 la1_data_in[1]
port 126 nsew signal input
rlabel metal3 s 0 32588 800 32828 6 la1_data_in[20]
port 127 nsew signal input
rlabel metal2 s 38630 49200 38742 50000 6 la1_data_in[21]
port 128 nsew signal input
rlabel metal3 s 39200 13548 40000 13788 6 la1_data_in[22]
port 129 nsew signal input
rlabel metal3 s 0 628 800 868 6 la1_data_in[23]
port 130 nsew signal input
rlabel metal2 s 12870 0 12982 800 6 la1_data_in[24]
port 131 nsew signal input
rlabel metal3 s 0 34628 800 34868 6 la1_data_in[25]
port 132 nsew signal input
rlabel metal3 s 39200 8108 40000 8348 6 la1_data_in[26]
port 133 nsew signal input
rlabel metal2 s 26394 0 26506 800 6 la1_data_in[27]
port 134 nsew signal input
rlabel metal3 s 0 29868 800 30108 6 la1_data_in[28]
port 135 nsew signal input
rlabel metal3 s 0 45508 800 45748 6 la1_data_in[29]
port 136 nsew signal input
rlabel metal2 s 10294 0 10406 800 6 la1_data_in[2]
port 137 nsew signal input
rlabel metal2 s 1278 0 1390 800 6 la1_data_in[30]
port 138 nsew signal input
rlabel metal2 s 34122 0 34234 800 6 la1_data_in[31]
port 139 nsew signal input
rlabel metal3 s 0 28508 800 28748 6 la1_data_in[3]
port 140 nsew signal input
rlabel metal2 s 32834 49200 32946 50000 6 la1_data_in[4]
port 141 nsew signal input
rlabel metal3 s 39200 27148 40000 27388 6 la1_data_in[5]
port 142 nsew signal input
rlabel metal2 s 12226 49200 12338 50000 6 la1_data_in[6]
port 143 nsew signal input
rlabel metal3 s 0 20348 800 20588 6 la1_data_in[7]
port 144 nsew signal input
rlabel metal2 s 12870 49200 12982 50000 6 la1_data_in[8]
port 145 nsew signal input
rlabel metal3 s 0 31228 800 31468 6 la1_data_in[9]
port 146 nsew signal input
rlabel metal2 s 7074 0 7186 800 6 la1_data_out[0]
port 147 nsew signal tristate
rlabel metal3 s 39200 15588 40000 15828 6 la1_data_out[10]
port 148 nsew signal tristate
rlabel metal2 s 20598 0 20710 800 6 la1_data_out[11]
port 149 nsew signal tristate
rlabel metal3 s 39200 46188 40000 46428 6 la1_data_out[12]
port 150 nsew signal tristate
rlabel metal3 s 0 49588 800 49828 6 la1_data_out[13]
port 151 nsew signal tristate
rlabel metal2 s 18666 49200 18778 50000 6 la1_data_out[14]
port 152 nsew signal tristate
rlabel metal3 s 0 1308 800 1548 6 la1_data_out[15]
port 153 nsew signal tristate
rlabel metal3 s 39200 20348 40000 20588 6 la1_data_out[16]
port 154 nsew signal tristate
rlabel metal3 s 39200 38028 40000 38268 6 la1_data_out[17]
port 155 nsew signal tristate
rlabel metal2 s -10 49200 102 50000 6 la1_data_out[18]
port 156 nsew signal tristate
rlabel metal3 s 39200 27828 40000 28068 6 la1_data_out[19]
port 157 nsew signal tristate
rlabel metal3 s 0 40748 800 40988 6 la1_data_out[1]
port 158 nsew signal tristate
rlabel metal3 s 0 9468 800 9708 6 la1_data_out[20]
port 159 nsew signal tristate
rlabel metal3 s 39200 44148 40000 44388 6 la1_data_out[21]
port 160 nsew signal tristate
rlabel metal2 s 22530 49200 22642 50000 6 la1_data_out[22]
port 161 nsew signal tristate
rlabel metal2 s 10938 0 11050 800 6 la1_data_out[23]
port 162 nsew signal tristate
rlabel metal3 s 39200 21708 40000 21948 6 la1_data_out[24]
port 163 nsew signal tristate
rlabel metal3 s 0 3348 800 3588 6 la1_data_out[25]
port 164 nsew signal tristate
rlabel metal3 s 39200 9468 40000 9708 6 la1_data_out[26]
port 165 nsew signal tristate
rlabel metal3 s 0 43468 800 43708 6 la1_data_out[27]
port 166 nsew signal tristate
rlabel metal3 s 39200 -52 40000 188 6 la1_data_out[28]
port 167 nsew signal tristate
rlabel metal2 s 5142 0 5254 800 6 la1_data_out[29]
port 168 nsew signal tristate
rlabel metal2 s 18666 0 18778 800 6 la1_data_out[2]
port 169 nsew signal tristate
rlabel metal3 s 39200 16948 40000 17188 6 la1_data_out[30]
port 170 nsew signal tristate
rlabel metal3 s 39200 48908 40000 49148 6 la1_data_out[31]
port 171 nsew signal tristate
rlabel metal3 s 0 8108 800 8348 6 la1_data_out[3]
port 172 nsew signal tristate
rlabel metal3 s 39200 1308 40000 1548 6 la1_data_out[4]
port 173 nsew signal tristate
rlabel metal2 s 3210 0 3322 800 6 la1_data_out[5]
port 174 nsew signal tristate
rlabel metal3 s 39200 23748 40000 23988 6 la1_data_out[6]
port 175 nsew signal tristate
rlabel metal2 s 634 0 746 800 6 la1_data_out[7]
port 176 nsew signal tristate
rlabel metal3 s 39200 38708 40000 38948 6 la1_data_out[8]
port 177 nsew signal tristate
rlabel metal2 s 37342 49200 37454 50000 6 la1_data_out[9]
port 178 nsew signal tristate
rlabel metal3 s 39200 4708 40000 4948 6 la1_oenb[0]
port 179 nsew signal input
rlabel metal2 s 35410 49200 35522 50000 6 la1_oenb[10]
port 180 nsew signal input
rlabel metal3 s 0 25108 800 25348 6 la1_oenb[11]
port 181 nsew signal input
rlabel metal3 s 0 26468 800 26708 6 la1_oenb[12]
port 182 nsew signal input
rlabel metal2 s 27038 0 27150 800 6 la1_oenb[13]
port 183 nsew signal input
rlabel metal2 s -10 0 102 800 6 la1_oenb[14]
port 184 nsew signal input
rlabel metal2 s 32190 0 32302 800 6 la1_oenb[15]
port 185 nsew signal input
rlabel metal3 s 0 31908 800 32148 6 la1_oenb[16]
port 186 nsew signal input
rlabel metal3 s 0 48228 800 48468 6 la1_oenb[17]
port 187 nsew signal input
rlabel metal2 s 14802 49200 14914 50000 6 la1_oenb[18]
port 188 nsew signal input
rlabel metal3 s 0 23748 800 23988 6 la1_oenb[19]
port 189 nsew signal input
rlabel metal2 s 7718 0 7830 800 6 la1_oenb[1]
port 190 nsew signal input
rlabel metal2 s 1922 0 2034 800 6 la1_oenb[20]
port 191 nsew signal input
rlabel metal2 s 23818 49200 23930 50000 6 la1_oenb[21]
port 192 nsew signal input
rlabel metal2 s 14158 49200 14270 50000 6 la1_oenb[22]
port 193 nsew signal input
rlabel metal2 s 21886 0 21998 800 6 la1_oenb[23]
port 194 nsew signal input
rlabel metal2 s 30258 49200 30370 50000 6 la1_oenb[24]
port 195 nsew signal input
rlabel metal3 s 39200 14228 40000 14468 6 la1_oenb[25]
port 196 nsew signal input
rlabel metal3 s 0 35308 800 35548 6 la1_oenb[26]
port 197 nsew signal input
rlabel metal3 s 39200 36668 40000 36908 6 la1_oenb[27]
port 198 nsew signal input
rlabel metal2 s 9006 0 9118 800 6 la1_oenb[28]
port 199 nsew signal input
rlabel metal2 s 16090 0 16202 800 6 la1_oenb[29]
port 200 nsew signal input
rlabel metal3 s 0 7428 800 7668 6 la1_oenb[2]
port 201 nsew signal input
rlabel metal3 s 39200 35988 40000 36228 6 la1_oenb[30]
port 202 nsew signal input
rlabel metal2 s 25106 0 25218 800 6 la1_oenb[31]
port 203 nsew signal input
rlabel metal2 s 26394 49200 26506 50000 6 la1_oenb[3]
port 204 nsew signal input
rlabel metal2 s 25750 49200 25862 50000 6 la1_oenb[4]
port 205 nsew signal input
rlabel metal3 s 0 44148 800 44388 6 la1_oenb[5]
port 206 nsew signal input
rlabel metal2 s 1278 49200 1390 50000 6 la1_oenb[6]
port 207 nsew signal input
rlabel metal2 s 30902 0 31014 800 6 la1_oenb[7]
port 208 nsew signal input
rlabel metal3 s 0 10828 800 11068 6 la1_oenb[8]
port 209 nsew signal input
rlabel metal3 s 0 38028 800 38268 6 la1_oenb[9]
port 210 nsew signal input
rlabel metal4 s 4208 2128 4528 47376 6 vccd1
port 211 nsew power input
rlabel metal4 s 34928 2128 35248 47376 6 vccd1
port 211 nsew power input
rlabel metal4 s 19568 2128 19888 47376 6 vssd1
port 212 nsew ground input
rlabel metal3 s 39200 26468 40000 26708 6 wb_clk_i
port 213 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 50000
<< end >>
